module sin_rom(
    clock,
    phase_in,
    sin_out,
);

// Input Ports
input clock;
input [11:0] phase_in;

// Output Ports
output [9:0] sin_out;

// Internal Ports
integer i;
reg [9:0] sine [0:4095];

initial begin
    sine[0]=0;
    sine[1]=1;
    sine[2]=3;
    sine[3]=4;
    sine[4]=6;
    sine[5]=7;
    sine[6]=9;
    sine[7]=10;
    sine[8]=12;
    sine[9]=14;
    sine[10]=15;
    sine[11]=17;
    sine[12]=18;
    sine[13]=20;
    sine[14]=21;
    sine[15]=23;
    sine[16]=25;
    sine[17]=26;
    sine[18]=28;
    sine[19]=29;
    sine[20]=31;
    sine[21]=32;
    sine[22]=34;
    sine[23]=36;
    sine[24]=37;
    sine[25]=39;
    sine[26]=40;
    sine[27]=42;
    sine[28]=43;
    sine[29]=45;
    sine[30]=47;
    sine[31]=48;
    sine[32]=50;
    sine[33]=51;
    sine[34]=53;
    sine[35]=54;
    sine[36]=56;
    sine[37]=58;
    sine[38]=59;
    sine[39]=61;
    sine[40]=62;
    sine[41]=64;
    sine[42]=65;
    sine[43]=67;
    sine[44]=69;
    sine[45]=70;
    sine[46]=72;
    sine[47]=73;
    sine[48]=75;
    sine[49]=76;
    sine[50]=78;
    sine[51]=80;
    sine[52]=81;
    sine[53]=83;
    sine[54]=84;
    sine[55]=86;
    sine[56]=87;
    sine[57]=89;
    sine[58]=90;
    sine[59]=92;
    sine[60]=94;
    sine[61]=95;
    sine[62]=97;
    sine[63]=98;
    sine[64]=100;
    sine[65]=101;
    sine[66]=103;
    sine[67]=105;
    sine[68]=106;
    sine[69]=108;
    sine[70]=109;
    sine[71]=111;
    sine[72]=112;
    sine[73]=114;
    sine[74]=115;
    sine[75]=117;
    sine[76]=119;
    sine[77]=120;
    sine[78]=122;
    sine[79]=123;
    sine[80]=125;
    sine[81]=126;
    sine[82]=128;
    sine[83]=130;
    sine[84]=131;
    sine[85]=133;
    sine[86]=134;
    sine[87]=136;
    sine[88]=137;
    sine[89]=139;
    sine[90]=140;
    sine[91]=142;
    sine[92]=144;
    sine[93]=145;
    sine[94]=147;
    sine[95]=148;
    sine[96]=150;
    sine[97]=151;
    sine[98]=153;
    sine[99]=154;
    sine[100]=156;
    sine[101]=158;
    sine[102]=159;
    sine[103]=161;
    sine[104]=162;
    sine[105]=164;
    sine[106]=165;
    sine[107]=167;
    sine[108]=168;
    sine[109]=170;
    sine[110]=171;
    sine[111]=173;
    sine[112]=175;
    sine[113]=176;
    sine[114]=178;
    sine[115]=179;
    sine[116]=181;
    sine[117]=182;
    sine[118]=184;
    sine[119]=185;
    sine[120]=187;
    sine[121]=188;
    sine[122]=190;
    sine[123]=192;
    sine[124]=193;
    sine[125]=195;
    sine[126]=196;
    sine[127]=198;
    sine[128]=199;
    sine[129]=201;
    sine[130]=202;
    sine[131]=204;
    sine[132]=205;
    sine[133]=207;
    sine[134]=209;
    sine[135]=210;
    sine[136]=212;
    sine[137]=213;
    sine[138]=215;
    sine[139]=216;
    sine[140]=218;
    sine[141]=219;
    sine[142]=221;
    sine[143]=222;
    sine[144]=224;
    sine[145]=225;
    sine[146]=227;
    sine[147]=228;
    sine[148]=230;
    sine[149]=232;
    sine[150]=233;
    sine[151]=235;
    sine[152]=236;
    sine[153]=238;
    sine[154]=239;
    sine[155]=241;
    sine[156]=242;
    sine[157]=244;
    sine[158]=245;
    sine[159]=247;
    sine[160]=248;
    sine[161]=250;
    sine[162]=251;
    sine[163]=253;
    sine[164]=254;
    sine[165]=256;
    sine[166]=257;
    sine[167]=259;
    sine[168]=260;
    sine[169]=262;
    sine[170]=264;
    sine[171]=265;
    sine[172]=267;
    sine[173]=268;
    sine[174]=270;
    sine[175]=271;
    sine[176]=273;
    sine[177]=274;
    sine[178]=276;
    sine[179]=277;
    sine[180]=279;
    sine[181]=280;
    sine[182]=282;
    sine[183]=283;
    sine[184]=285;
    sine[185]=286;
    sine[186]=288;
    sine[187]=289;
    sine[188]=291;
    sine[189]=292;
    sine[190]=294;
    sine[191]=295;
    sine[192]=297;
    sine[193]=298;
    sine[194]=300;
    sine[195]=301;
    sine[196]=303;
    sine[197]=304;
    sine[198]=306;
    sine[199]=307;
    sine[200]=309;
    sine[201]=310;
    sine[202]=312;
    sine[203]=313;
    sine[204]=315;
    sine[205]=316;
    sine[206]=318;
    sine[207]=319;
    sine[208]=321;
    sine[209]=322;
    sine[210]=324;
    sine[211]=325;
    sine[212]=327;
    sine[213]=328;
    sine[214]=330;
    sine[215]=331;
    sine[216]=333;
    sine[217]=334;
    sine[218]=336;
    sine[219]=337;
    sine[220]=339;
    sine[221]=340;
    sine[222]=342;
    sine[223]=343;
    sine[224]=344;
    sine[225]=346;
    sine[226]=347;
    sine[227]=349;
    sine[228]=350;
    sine[229]=352;
    sine[230]=353;
    sine[231]=355;
    sine[232]=356;
    sine[233]=358;
    sine[234]=359;
    sine[235]=361;
    sine[236]=362;
    sine[237]=364;
    sine[238]=365;
    sine[239]=367;
    sine[240]=368;
    sine[241]=369;
    sine[242]=371;
    sine[243]=372;
    sine[244]=374;
    sine[245]=375;
    sine[246]=377;
    sine[247]=378;
    sine[248]=380;
    sine[249]=381;
    sine[250]=383;
    sine[251]=384;
    sine[252]=386;
    sine[253]=387;
    sine[254]=388;
    sine[255]=390;
    sine[256]=391;
    sine[257]=393;
    sine[258]=394;
    sine[259]=396;
    sine[260]=397;
    sine[261]=399;
    sine[262]=400;
    sine[263]=402;
    sine[264]=403;
    sine[265]=404;
    sine[266]=406;
    sine[267]=407;
    sine[268]=409;
    sine[269]=410;
    sine[270]=412;
    sine[271]=413;
    sine[272]=414;
    sine[273]=416;
    sine[274]=417;
    sine[275]=419;
    sine[276]=420;
    sine[277]=422;
    sine[278]=423;
    sine[279]=424;
    sine[280]=426;
    sine[281]=427;
    sine[282]=429;
    sine[283]=430;
    sine[284]=432;
    sine[285]=433;
    sine[286]=434;
    sine[287]=436;
    sine[288]=437;
    sine[289]=439;
    sine[290]=440;
    sine[291]=442;
    sine[292]=443;
    sine[293]=444;
    sine[294]=446;
    sine[295]=447;
    sine[296]=449;
    sine[297]=450;
    sine[298]=451;
    sine[299]=453;
    sine[300]=454;
    sine[301]=456;
    sine[302]=457;
    sine[303]=458;
    sine[304]=460;
    sine[305]=461;
    sine[306]=463;
    sine[307]=464;
    sine[308]=466;
    sine[309]=467;
    sine[310]=468;
    sine[311]=470;
    sine[312]=471;
    sine[313]=472;
    sine[314]=474;
    sine[315]=475;
    sine[316]=477;
    sine[317]=478;
    sine[318]=479;
    sine[319]=481;
    sine[320]=482;
    sine[321]=484;
    sine[322]=485;
    sine[323]=486;
    sine[324]=488;
    sine[325]=489;
    sine[326]=491;
    sine[327]=492;
    sine[328]=493;
    sine[329]=495;
    sine[330]=496;
    sine[331]=497;
    sine[332]=499;
    sine[333]=500;
    sine[334]=501;
    sine[335]=503;
    sine[336]=504;
    sine[337]=506;
    sine[338]=507;
    sine[339]=508;
    sine[340]=510;
    sine[341]=511;
    sine[342]=512;
    sine[343]=514;
    sine[344]=515;
    sine[345]=516;
    sine[346]=518;
    sine[347]=519;
    sine[348]=521;
    sine[349]=522;
    sine[350]=523;
    sine[351]=525;
    sine[352]=526;
    sine[353]=527;
    sine[354]=529;
    sine[355]=530;
    sine[356]=531;
    sine[357]=533;
    sine[358]=534;
    sine[359]=535;
    sine[360]=537;
    sine[361]=538;
    sine[362]=539;
    sine[363]=541;
    sine[364]=542;
    sine[365]=543;
    sine[366]=545;
    sine[367]=546;
    sine[368]=547;
    sine[369]=549;
    sine[370]=550;
    sine[371]=551;
    sine[372]=553;
    sine[373]=554;
    sine[374]=555;
    sine[375]=557;
    sine[376]=558;
    sine[377]=559;
    sine[378]=561;
    sine[379]=562;
    sine[380]=563;
    sine[381]=564;
    sine[382]=566;
    sine[383]=567;
    sine[384]=568;
    sine[385]=570;
    sine[386]=571;
    sine[387]=572;
    sine[388]=574;
    sine[389]=575;
    sine[390]=576;
    sine[391]=578;
    sine[392]=579;
    sine[393]=580;
    sine[394]=581;
    sine[395]=583;
    sine[396]=584;
    sine[397]=585;
    sine[398]=587;
    sine[399]=588;
    sine[400]=589;
    sine[401]=590;
    sine[402]=592;
    sine[403]=593;
    sine[404]=594;
    sine[405]=596;
    sine[406]=597;
    sine[407]=598;
    sine[408]=599;
    sine[409]=601;
    sine[410]=602;
    sine[411]=603;
    sine[412]=604;
    sine[413]=606;
    sine[414]=607;
    sine[415]=608;
    sine[416]=609;
    sine[417]=611;
    sine[418]=612;
    sine[419]=613;
    sine[420]=615;
    sine[421]=616;
    sine[422]=617;
    sine[423]=618;
    sine[424]=620;
    sine[425]=621;
    sine[426]=622;
    sine[427]=623;
    sine[428]=625;
    sine[429]=626;
    sine[430]=627;
    sine[431]=628;
    sine[432]=629;
    sine[433]=631;
    sine[434]=632;
    sine[435]=633;
    sine[436]=634;
    sine[437]=636;
    sine[438]=637;
    sine[439]=638;
    sine[440]=639;
    sine[441]=641;
    sine[442]=642;
    sine[443]=643;
    sine[444]=644;
    sine[445]=645;
    sine[446]=647;
    sine[447]=648;
    sine[448]=649;
    sine[449]=650;
    sine[450]=652;
    sine[451]=653;
    sine[452]=654;
    sine[453]=655;
    sine[454]=656;
    sine[455]=658;
    sine[456]=659;
    sine[457]=660;
    sine[458]=661;
    sine[459]=662;
    sine[460]=664;
    sine[461]=665;
    sine[462]=666;
    sine[463]=667;
    sine[464]=668;
    sine[465]=670;
    sine[466]=671;
    sine[467]=672;
    sine[468]=673;
    sine[469]=674;
    sine[470]=675;
    sine[471]=677;
    sine[472]=678;
    sine[473]=679;
    sine[474]=680;
    sine[475]=681;
    sine[476]=683;
    sine[477]=684;
    sine[478]=685;
    sine[479]=686;
    sine[480]=687;
    sine[481]=688;
    sine[482]=690;
    sine[483]=691;
    sine[484]=692;
    sine[485]=693;
    sine[486]=694;
    sine[487]=695;
    sine[488]=696;
    sine[489]=698;
    sine[490]=699;
    sine[491]=700;
    sine[492]=701;
    sine[493]=702;
    sine[494]=703;
    sine[495]=704;
    sine[496]=706;
    sine[497]=707;
    sine[498]=708;
    sine[499]=709;
    sine[500]=710;
    sine[501]=711;
    sine[502]=712;
    sine[503]=714;
    sine[504]=715;
    sine[505]=716;
    sine[506]=717;
    sine[507]=718;
    sine[508]=719;
    sine[509]=720;
    sine[510]=721;
    sine[511]=722;
    sine[512]=724;
    sine[513]=725;
    sine[514]=726;
    sine[515]=727;
    sine[516]=728;
    sine[517]=729;
    sine[518]=730;
    sine[519]=731;
    sine[520]=732;
    sine[521]=734;
    sine[522]=735;
    sine[523]=736;
    sine[524]=737;
    sine[525]=738;
    sine[526]=739;
    sine[527]=740;
    sine[528]=741;
    sine[529]=742;
    sine[530]=743;
    sine[531]=744;
    sine[532]=745;
    sine[533]=747;
    sine[534]=748;
    sine[535]=749;
    sine[536]=750;
    sine[537]=751;
    sine[538]=752;
    sine[539]=753;
    sine[540]=754;
    sine[541]=755;
    sine[542]=756;
    sine[543]=757;
    sine[544]=758;
    sine[545]=759;
    sine[546]=760;
    sine[547]=761;
    sine[548]=762;
    sine[549]=763;
    sine[550]=765;
    sine[551]=766;
    sine[552]=767;
    sine[553]=768;
    sine[554]=769;
    sine[555]=770;
    sine[556]=771;
    sine[557]=772;
    sine[558]=773;
    sine[559]=774;
    sine[560]=775;
    sine[561]=776;
    sine[562]=777;
    sine[563]=778;
    sine[564]=779;
    sine[565]=780;
    sine[566]=781;
    sine[567]=782;
    sine[568]=783;
    sine[569]=784;
    sine[570]=785;
    sine[571]=786;
    sine[572]=787;
    sine[573]=788;
    sine[574]=789;
    sine[575]=790;
    sine[576]=791;
    sine[577]=792;
    sine[578]=793;
    sine[579]=794;
    sine[580]=795;
    sine[581]=796;
    sine[582]=797;
    sine[583]=798;
    sine[584]=799;
    sine[585]=800;
    sine[586]=801;
    sine[587]=802;
    sine[588]=803;
    sine[589]=804;
    sine[590]=805;
    sine[591]=806;
    sine[592]=807;
    sine[593]=808;
    sine[594]=809;
    sine[595]=810;
    sine[596]=811;
    sine[597]=812;
    sine[598]=813;
    sine[599]=813;
    sine[600]=814;
    sine[601]=815;
    sine[602]=816;
    sine[603]=817;
    sine[604]=818;
    sine[605]=819;
    sine[606]=820;
    sine[607]=821;
    sine[608]=822;
    sine[609]=823;
    sine[610]=824;
    sine[611]=825;
    sine[612]=826;
    sine[613]=827;
    sine[614]=828;
    sine[615]=828;
    sine[616]=829;
    sine[617]=830;
    sine[618]=831;
    sine[619]=832;
    sine[620]=833;
    sine[621]=834;
    sine[622]=835;
    sine[623]=836;
    sine[624]=837;
    sine[625]=838;
    sine[626]=839;
    sine[627]=839;
    sine[628]=840;
    sine[629]=841;
    sine[630]=842;
    sine[631]=843;
    sine[632]=844;
    sine[633]=845;
    sine[634]=846;
    sine[635]=847;
    sine[636]=847;
    sine[637]=848;
    sine[638]=849;
    sine[639]=850;
    sine[640]=851;
    sine[641]=852;
    sine[642]=853;
    sine[643]=854;
    sine[644]=854;
    sine[645]=855;
    sine[646]=856;
    sine[647]=857;
    sine[648]=858;
    sine[649]=859;
    sine[650]=860;
    sine[651]=860;
    sine[652]=861;
    sine[653]=862;
    sine[654]=863;
    sine[655]=864;
    sine[656]=865;
    sine[657]=865;
    sine[658]=866;
    sine[659]=867;
    sine[660]=868;
    sine[661]=869;
    sine[662]=870;
    sine[663]=870;
    sine[664]=871;
    sine[665]=872;
    sine[666]=873;
    sine[667]=874;
    sine[668]=875;
    sine[669]=875;
    sine[670]=876;
    sine[671]=877;
    sine[672]=878;
    sine[673]=879;
    sine[674]=879;
    sine[675]=880;
    sine[676]=881;
    sine[677]=882;
    sine[678]=883;
    sine[679]=883;
    sine[680]=884;
    sine[681]=885;
    sine[682]=886;
    sine[683]=887;
    sine[684]=887;
    sine[685]=888;
    sine[686]=889;
    sine[687]=890;
    sine[688]=890;
    sine[689]=891;
    sine[690]=892;
    sine[691]=893;
    sine[692]=894;
    sine[693]=894;
    sine[694]=895;
    sine[695]=896;
    sine[696]=897;
    sine[697]=897;
    sine[698]=898;
    sine[699]=899;
    sine[700]=900;
    sine[701]=900;
    sine[702]=901;
    sine[703]=902;
    sine[704]=903;
    sine[705]=903;
    sine[706]=904;
    sine[707]=905;
    sine[708]=906;
    sine[709]=906;
    sine[710]=907;
    sine[711]=908;
    sine[712]=908;
    sine[713]=909;
    sine[714]=910;
    sine[715]=911;
    sine[716]=911;
    sine[717]=912;
    sine[718]=913;
    sine[719]=913;
    sine[720]=914;
    sine[721]=915;
    sine[722]=916;
    sine[723]=916;
    sine[724]=917;
    sine[725]=918;
    sine[726]=918;
    sine[727]=919;
    sine[728]=920;
    sine[729]=920;
    sine[730]=921;
    sine[731]=922;
    sine[732]=922;
    sine[733]=923;
    sine[734]=924;
    sine[735]=925;
    sine[736]=925;
    sine[737]=926;
    sine[738]=927;
    sine[739]=927;
    sine[740]=928;
    sine[741]=929;
    sine[742]=929;
    sine[743]=930;
    sine[744]=930;
    sine[745]=931;
    sine[746]=932;
    sine[747]=932;
    sine[748]=933;
    sine[749]=934;
    sine[750]=934;
    sine[751]=935;
    sine[752]=936;
    sine[753]=936;
    sine[754]=937;
    sine[755]=938;
    sine[756]=938;
    sine[757]=939;
    sine[758]=939;
    sine[759]=940;
    sine[760]=941;
    sine[761]=941;
    sine[762]=942;
    sine[763]=943;
    sine[764]=943;
    sine[765]=944;
    sine[766]=944;
    sine[767]=945;
    sine[768]=946;
    sine[769]=946;
    sine[770]=947;
    sine[771]=947;
    sine[772]=948;
    sine[773]=949;
    sine[774]=949;
    sine[775]=950;
    sine[776]=950;
    sine[777]=951;
    sine[778]=951;
    sine[779]=952;
    sine[780]=953;
    sine[781]=953;
    sine[782]=954;
    sine[783]=954;
    sine[784]=955;
    sine[785]=955;
    sine[786]=956;
    sine[787]=957;
    sine[788]=957;
    sine[789]=958;
    sine[790]=958;
    sine[791]=959;
    sine[792]=959;
    sine[793]=960;
    sine[794]=960;
    sine[795]=961;
    sine[796]=962;
    sine[797]=962;
    sine[798]=963;
    sine[799]=963;
    sine[800]=964;
    sine[801]=964;
    sine[802]=965;
    sine[803]=965;
    sine[804]=966;
    sine[805]=966;
    sine[806]=967;
    sine[807]=967;
    sine[808]=968;
    sine[809]=968;
    sine[810]=969;
    sine[811]=969;
    sine[812]=970;
    sine[813]=970;
    sine[814]=971;
    sine[815]=971;
    sine[816]=972;
    sine[817]=972;
    sine[818]=973;
    sine[819]=973;
    sine[820]=974;
    sine[821]=974;
    sine[822]=975;
    sine[823]=975;
    sine[824]=976;
    sine[825]=976;
    sine[826]=977;
    sine[827]=977;
    sine[828]=978;
    sine[829]=978;
    sine[830]=978;
    sine[831]=979;
    sine[832]=979;
    sine[833]=980;
    sine[834]=980;
    sine[835]=981;
    sine[836]=981;
    sine[837]=982;
    sine[838]=982;
    sine[839]=983;
    sine[840]=983;
    sine[841]=983;
    sine[842]=984;
    sine[843]=984;
    sine[844]=985;
    sine[845]=985;
    sine[846]=986;
    sine[847]=986;
    sine[848]=986;
    sine[849]=987;
    sine[850]=987;
    sine[851]=988;
    sine[852]=988;
    sine[853]=988;
    sine[854]=989;
    sine[855]=989;
    sine[856]=990;
    sine[857]=990;
    sine[858]=990;
    sine[859]=991;
    sine[860]=991;
    sine[861]=992;
    sine[862]=992;
    sine[863]=992;
    sine[864]=993;
    sine[865]=993;
    sine[866]=994;
    sine[867]=994;
    sine[868]=994;
    sine[869]=995;
    sine[870]=995;
    sine[871]=995;
    sine[872]=996;
    sine[873]=996;
    sine[874]=997;
    sine[875]=997;
    sine[876]=997;
    sine[877]=998;
    sine[878]=998;
    sine[879]=998;
    sine[880]=999;
    sine[881]=999;
    sine[882]=999;
    sine[883]=1000;
    sine[884]=1000;
    sine[885]=1000;
    sine[886]=1001;
    sine[887]=1001;
    sine[888]=1001;
    sine[889]=1002;
    sine[890]=1002;
    sine[891]=1002;
    sine[892]=1003;
    sine[893]=1003;
    sine[894]=1003;
    sine[895]=1004;
    sine[896]=1004;
    sine[897]=1004;
    sine[898]=1004;
    sine[899]=1005;
    sine[900]=1005;
    sine[901]=1005;
    sine[902]=1006;
    sine[903]=1006;
    sine[904]=1006;
    sine[905]=1006;
    sine[906]=1007;
    sine[907]=1007;
    sine[908]=1007;
    sine[909]=1008;
    sine[910]=1008;
    sine[911]=1008;
    sine[912]=1008;
    sine[913]=1009;
    sine[914]=1009;
    sine[915]=1009;
    sine[916]=1009;
    sine[917]=1010;
    sine[918]=1010;
    sine[919]=1010;
    sine[920]=1010;
    sine[921]=1011;
    sine[922]=1011;
    sine[923]=1011;
    sine[924]=1011;
    sine[925]=1012;
    sine[926]=1012;
    sine[927]=1012;
    sine[928]=1012;
    sine[929]=1013;
    sine[930]=1013;
    sine[931]=1013;
    sine[932]=1013;
    sine[933]=1014;
    sine[934]=1014;
    sine[935]=1014;
    sine[936]=1014;
    sine[937]=1014;
    sine[938]=1015;
    sine[939]=1015;
    sine[940]=1015;
    sine[941]=1015;
    sine[942]=1015;
    sine[943]=1016;
    sine[944]=1016;
    sine[945]=1016;
    sine[946]=1016;
    sine[947]=1016;
    sine[948]=1017;
    sine[949]=1017;
    sine[950]=1017;
    sine[951]=1017;
    sine[952]=1017;
    sine[953]=1017;
    sine[954]=1018;
    sine[955]=1018;
    sine[956]=1018;
    sine[957]=1018;
    sine[958]=1018;
    sine[959]=1018;
    sine[960]=1019;
    sine[961]=1019;
    sine[962]=1019;
    sine[963]=1019;
    sine[964]=1019;
    sine[965]=1019;
    sine[966]=1019;
    sine[967]=1020;
    sine[968]=1020;
    sine[969]=1020;
    sine[970]=1020;
    sine[971]=1020;
    sine[972]=1020;
    sine[973]=1020;
    sine[974]=1020;
    sine[975]=1021;
    sine[976]=1021;
    sine[977]=1021;
    sine[978]=1021;
    sine[979]=1021;
    sine[980]=1021;
    sine[981]=1021;
    sine[982]=1021;
    sine[983]=1021;
    sine[984]=1022;
    sine[985]=1022;
    sine[986]=1022;
    sine[987]=1022;
    sine[988]=1022;
    sine[989]=1022;
    sine[990]=1022;
    sine[991]=1022;
    sine[992]=1022;
    sine[993]=1022;
    sine[994]=1022;
    sine[995]=1022;
    sine[996]=1023;
    sine[997]=1023;
    sine[998]=1023;
    sine[999]=1023;
    sine[1000]=1023;
    sine[1001]=1023;
    sine[1002]=1023;
    sine[1003]=1023;
    sine[1004]=1023;
    sine[1005]=1023;
    sine[1006]=1023;
    sine[1007]=1023;
    sine[1008]=1023;
    sine[1009]=1023;
    sine[1010]=1023;
    sine[1011]=1023;
    sine[1012]=1023;
    sine[1013]=1023;
    sine[1014]=1023;
    sine[1015]=1023;
    sine[1016]=1023;
    sine[1017]=1023;
    sine[1018]=1023;
    sine[1019]=1023;
    sine[1020]=1023;
    sine[1021]=1023;
    sine[1022]=1023;
    sine[1023]=1023;
    sine[1024]=1024;
    sine[1025]=1023;
    sine[1026]=1023;
    sine[1027]=1023;
    sine[1028]=1023;
    sine[1029]=1023;
    sine[1030]=1023;
    sine[1031]=1023;
    sine[1032]=1023;
    sine[1033]=1023;
    sine[1034]=1023;
    sine[1035]=1023;
    sine[1036]=1023;
    sine[1037]=1023;
    sine[1038]=1023;
    sine[1039]=1023;
    sine[1040]=1023;
    sine[1041]=1023;
    sine[1042]=1023;
    sine[1043]=1023;
    sine[1044]=1023;
    sine[1045]=1023;
    sine[1046]=1023;
    sine[1047]=1023;
    sine[1048]=1023;
    sine[1049]=1023;
    sine[1050]=1023;
    sine[1051]=1023;
    sine[1052]=1023;
    sine[1053]=1022;
    sine[1054]=1022;
    sine[1055]=1022;
    sine[1056]=1022;
    sine[1057]=1022;
    sine[1058]=1022;
    sine[1059]=1022;
    sine[1060]=1022;
    sine[1061]=1022;
    sine[1062]=1022;
    sine[1063]=1022;
    sine[1064]=1022;
    sine[1065]=1021;
    sine[1066]=1021;
    sine[1067]=1021;
    sine[1068]=1021;
    sine[1069]=1021;
    sine[1070]=1021;
    sine[1071]=1021;
    sine[1072]=1021;
    sine[1073]=1021;
    sine[1074]=1020;
    sine[1075]=1020;
    sine[1076]=1020;
    sine[1077]=1020;
    sine[1078]=1020;
    sine[1079]=1020;
    sine[1080]=1020;
    sine[1081]=1020;
    sine[1082]=1019;
    sine[1083]=1019;
    sine[1084]=1019;
    sine[1085]=1019;
    sine[1086]=1019;
    sine[1087]=1019;
    sine[1088]=1019;
    sine[1089]=1018;
    sine[1090]=1018;
    sine[1091]=1018;
    sine[1092]=1018;
    sine[1093]=1018;
    sine[1094]=1018;
    sine[1095]=1017;
    sine[1096]=1017;
    sine[1097]=1017;
    sine[1098]=1017;
    sine[1099]=1017;
    sine[1100]=1017;
    sine[1101]=1016;
    sine[1102]=1016;
    sine[1103]=1016;
    sine[1104]=1016;
    sine[1105]=1016;
    sine[1106]=1015;
    sine[1107]=1015;
    sine[1108]=1015;
    sine[1109]=1015;
    sine[1110]=1015;
    sine[1111]=1014;
    sine[1112]=1014;
    sine[1113]=1014;
    sine[1114]=1014;
    sine[1115]=1014;
    sine[1116]=1013;
    sine[1117]=1013;
    sine[1118]=1013;
    sine[1119]=1013;
    sine[1120]=1012;
    sine[1121]=1012;
    sine[1122]=1012;
    sine[1123]=1012;
    sine[1124]=1011;
    sine[1125]=1011;
    sine[1126]=1011;
    sine[1127]=1011;
    sine[1128]=1010;
    sine[1129]=1010;
    sine[1130]=1010;
    sine[1131]=1010;
    sine[1132]=1009;
    sine[1133]=1009;
    sine[1134]=1009;
    sine[1135]=1009;
    sine[1136]=1008;
    sine[1137]=1008;
    sine[1138]=1008;
    sine[1139]=1008;
    sine[1140]=1007;
    sine[1141]=1007;
    sine[1142]=1007;
    sine[1143]=1006;
    sine[1144]=1006;
    sine[1145]=1006;
    sine[1146]=1006;
    sine[1147]=1005;
    sine[1148]=1005;
    sine[1149]=1005;
    sine[1150]=1004;
    sine[1151]=1004;
    sine[1152]=1004;
    sine[1153]=1004;
    sine[1154]=1003;
    sine[1155]=1003;
    sine[1156]=1003;
    sine[1157]=1002;
    sine[1158]=1002;
    sine[1159]=1002;
    sine[1160]=1001;
    sine[1161]=1001;
    sine[1162]=1001;
    sine[1163]=1000;
    sine[1164]=1000;
    sine[1165]=1000;
    sine[1166]=999;
    sine[1167]=999;
    sine[1168]=999;
    sine[1169]=998;
    sine[1170]=998;
    sine[1171]=998;
    sine[1172]=997;
    sine[1173]=997;
    sine[1174]=997;
    sine[1175]=996;
    sine[1176]=996;
    sine[1177]=995;
    sine[1178]=995;
    sine[1179]=995;
    sine[1180]=994;
    sine[1181]=994;
    sine[1182]=994;
    sine[1183]=993;
    sine[1184]=993;
    sine[1185]=992;
    sine[1186]=992;
    sine[1187]=992;
    sine[1188]=991;
    sine[1189]=991;
    sine[1190]=990;
    sine[1191]=990;
    sine[1192]=990;
    sine[1193]=989;
    sine[1194]=989;
    sine[1195]=988;
    sine[1196]=988;
    sine[1197]=988;
    sine[1198]=987;
    sine[1199]=987;
    sine[1200]=986;
    sine[1201]=986;
    sine[1202]=986;
    sine[1203]=985;
    sine[1204]=985;
    sine[1205]=984;
    sine[1206]=984;
    sine[1207]=983;
    sine[1208]=983;
    sine[1209]=983;
    sine[1210]=982;
    sine[1211]=982;
    sine[1212]=981;
    sine[1213]=981;
    sine[1214]=980;
    sine[1215]=980;
    sine[1216]=979;
    sine[1217]=979;
    sine[1218]=978;
    sine[1219]=978;
    sine[1220]=978;
    sine[1221]=977;
    sine[1222]=977;
    sine[1223]=976;
    sine[1224]=976;
    sine[1225]=975;
    sine[1226]=975;
    sine[1227]=974;
    sine[1228]=974;
    sine[1229]=973;
    sine[1230]=973;
    sine[1231]=972;
    sine[1232]=972;
    sine[1233]=971;
    sine[1234]=971;
    sine[1235]=970;
    sine[1236]=970;
    sine[1237]=969;
    sine[1238]=969;
    sine[1239]=968;
    sine[1240]=968;
    sine[1241]=967;
    sine[1242]=967;
    sine[1243]=966;
    sine[1244]=966;
    sine[1245]=965;
    sine[1246]=965;
    sine[1247]=964;
    sine[1248]=964;
    sine[1249]=963;
    sine[1250]=963;
    sine[1251]=962;
    sine[1252]=962;
    sine[1253]=961;
    sine[1254]=960;
    sine[1255]=960;
    sine[1256]=959;
    sine[1257]=959;
    sine[1258]=958;
    sine[1259]=958;
    sine[1260]=957;
    sine[1261]=957;
    sine[1262]=956;
    sine[1263]=955;
    sine[1264]=955;
    sine[1265]=954;
    sine[1266]=954;
    sine[1267]=953;
    sine[1268]=953;
    sine[1269]=952;
    sine[1270]=951;
    sine[1271]=951;
    sine[1272]=950;
    sine[1273]=950;
    sine[1274]=949;
    sine[1275]=949;
    sine[1276]=948;
    sine[1277]=947;
    sine[1278]=947;
    sine[1279]=946;
    sine[1280]=946;
    sine[1281]=945;
    sine[1282]=944;
    sine[1283]=944;
    sine[1284]=943;
    sine[1285]=943;
    sine[1286]=942;
    sine[1287]=941;
    sine[1288]=941;
    sine[1289]=940;
    sine[1290]=939;
    sine[1291]=939;
    sine[1292]=938;
    sine[1293]=938;
    sine[1294]=937;
    sine[1295]=936;
    sine[1296]=936;
    sine[1297]=935;
    sine[1298]=934;
    sine[1299]=934;
    sine[1300]=933;
    sine[1301]=932;
    sine[1302]=932;
    sine[1303]=931;
    sine[1304]=930;
    sine[1305]=930;
    sine[1306]=929;
    sine[1307]=929;
    sine[1308]=928;
    sine[1309]=927;
    sine[1310]=927;
    sine[1311]=926;
    sine[1312]=925;
    sine[1313]=925;
    sine[1314]=924;
    sine[1315]=923;
    sine[1316]=922;
    sine[1317]=922;
    sine[1318]=921;
    sine[1319]=920;
    sine[1320]=920;
    sine[1321]=919;
    sine[1322]=918;
    sine[1323]=918;
    sine[1324]=917;
    sine[1325]=916;
    sine[1326]=916;
    sine[1327]=915;
    sine[1328]=914;
    sine[1329]=913;
    sine[1330]=913;
    sine[1331]=912;
    sine[1332]=911;
    sine[1333]=911;
    sine[1334]=910;
    sine[1335]=909;
    sine[1336]=908;
    sine[1337]=908;
    sine[1338]=907;
    sine[1339]=906;
    sine[1340]=906;
    sine[1341]=905;
    sine[1342]=904;
    sine[1343]=903;
    sine[1344]=903;
    sine[1345]=902;
    sine[1346]=901;
    sine[1347]=900;
    sine[1348]=900;
    sine[1349]=899;
    sine[1350]=898;
    sine[1351]=897;
    sine[1352]=897;
    sine[1353]=896;
    sine[1354]=895;
    sine[1355]=894;
    sine[1356]=894;
    sine[1357]=893;
    sine[1358]=892;
    sine[1359]=891;
    sine[1360]=890;
    sine[1361]=890;
    sine[1362]=889;
    sine[1363]=888;
    sine[1364]=887;
    sine[1365]=887;
    sine[1366]=886;
    sine[1367]=885;
    sine[1368]=884;
    sine[1369]=883;
    sine[1370]=883;
    sine[1371]=882;
    sine[1372]=881;
    sine[1373]=880;
    sine[1374]=879;
    sine[1375]=879;
    sine[1376]=878;
    sine[1377]=877;
    sine[1378]=876;
    sine[1379]=875;
    sine[1380]=875;
    sine[1381]=874;
    sine[1382]=873;
    sine[1383]=872;
    sine[1384]=871;
    sine[1385]=870;
    sine[1386]=870;
    sine[1387]=869;
    sine[1388]=868;
    sine[1389]=867;
    sine[1390]=866;
    sine[1391]=865;
    sine[1392]=865;
    sine[1393]=864;
    sine[1394]=863;
    sine[1395]=862;
    sine[1396]=861;
    sine[1397]=860;
    sine[1398]=860;
    sine[1399]=859;
    sine[1400]=858;
    sine[1401]=857;
    sine[1402]=856;
    sine[1403]=855;
    sine[1404]=854;
    sine[1405]=854;
    sine[1406]=853;
    sine[1407]=852;
    sine[1408]=851;
    sine[1409]=850;
    sine[1410]=849;
    sine[1411]=848;
    sine[1412]=847;
    sine[1413]=847;
    sine[1414]=846;
    sine[1415]=845;
    sine[1416]=844;
    sine[1417]=843;
    sine[1418]=842;
    sine[1419]=841;
    sine[1420]=840;
    sine[1421]=839;
    sine[1422]=839;
    sine[1423]=838;
    sine[1424]=837;
    sine[1425]=836;
    sine[1426]=835;
    sine[1427]=834;
    sine[1428]=833;
    sine[1429]=832;
    sine[1430]=831;
    sine[1431]=830;
    sine[1432]=829;
    sine[1433]=828;
    sine[1434]=828;
    sine[1435]=827;
    sine[1436]=826;
    sine[1437]=825;
    sine[1438]=824;
    sine[1439]=823;
    sine[1440]=822;
    sine[1441]=821;
    sine[1442]=820;
    sine[1443]=819;
    sine[1444]=818;
    sine[1445]=817;
    sine[1446]=816;
    sine[1447]=815;
    sine[1448]=814;
    sine[1449]=813;
    sine[1450]=813;
    sine[1451]=812;
    sine[1452]=811;
    sine[1453]=810;
    sine[1454]=809;
    sine[1455]=808;
    sine[1456]=807;
    sine[1457]=806;
    sine[1458]=805;
    sine[1459]=804;
    sine[1460]=803;
    sine[1461]=802;
    sine[1462]=801;
    sine[1463]=800;
    sine[1464]=799;
    sine[1465]=798;
    sine[1466]=797;
    sine[1467]=796;
    sine[1468]=795;
    sine[1469]=794;
    sine[1470]=793;
    sine[1471]=792;
    sine[1472]=791;
    sine[1473]=790;
    sine[1474]=789;
    sine[1475]=788;
    sine[1476]=787;
    sine[1477]=786;
    sine[1478]=785;
    sine[1479]=784;
    sine[1480]=783;
    sine[1481]=782;
    sine[1482]=781;
    sine[1483]=780;
    sine[1484]=779;
    sine[1485]=778;
    sine[1486]=777;
    sine[1487]=776;
    sine[1488]=775;
    sine[1489]=774;
    sine[1490]=773;
    sine[1491]=772;
    sine[1492]=771;
    sine[1493]=770;
    sine[1494]=769;
    sine[1495]=768;
    sine[1496]=767;
    sine[1497]=766;
    sine[1498]=765;
    sine[1499]=763;
    sine[1500]=762;
    sine[1501]=761;
    sine[1502]=760;
    sine[1503]=759;
    sine[1504]=758;
    sine[1505]=757;
    sine[1506]=756;
    sine[1507]=755;
    sine[1508]=754;
    sine[1509]=753;
    sine[1510]=752;
    sine[1511]=751;
    sine[1512]=750;
    sine[1513]=749;
    sine[1514]=748;
    sine[1515]=747;
    sine[1516]=745;
    sine[1517]=744;
    sine[1518]=743;
    sine[1519]=742;
    sine[1520]=741;
    sine[1521]=740;
    sine[1522]=739;
    sine[1523]=738;
    sine[1524]=737;
    sine[1525]=736;
    sine[1526]=735;
    sine[1527]=734;
    sine[1528]=732;
    sine[1529]=731;
    sine[1530]=730;
    sine[1531]=729;
    sine[1532]=728;
    sine[1533]=727;
    sine[1534]=726;
    sine[1535]=725;
    sine[1536]=724;
    sine[1537]=722;
    sine[1538]=721;
    sine[1539]=720;
    sine[1540]=719;
    sine[1541]=718;
    sine[1542]=717;
    sine[1543]=716;
    sine[1544]=715;
    sine[1545]=714;
    sine[1546]=712;
    sine[1547]=711;
    sine[1548]=710;
    sine[1549]=709;
    sine[1550]=708;
    sine[1551]=707;
    sine[1552]=706;
    sine[1553]=704;
    sine[1554]=703;
    sine[1555]=702;
    sine[1556]=701;
    sine[1557]=700;
    sine[1558]=699;
    sine[1559]=698;
    sine[1560]=696;
    sine[1561]=695;
    sine[1562]=694;
    sine[1563]=693;
    sine[1564]=692;
    sine[1565]=691;
    sine[1566]=690;
    sine[1567]=688;
    sine[1568]=687;
    sine[1569]=686;
    sine[1570]=685;
    sine[1571]=684;
    sine[1572]=683;
    sine[1573]=681;
    sine[1574]=680;
    sine[1575]=679;
    sine[1576]=678;
    sine[1577]=677;
    sine[1578]=675;
    sine[1579]=674;
    sine[1580]=673;
    sine[1581]=672;
    sine[1582]=671;
    sine[1583]=670;
    sine[1584]=668;
    sine[1585]=667;
    sine[1586]=666;
    sine[1587]=665;
    sine[1588]=664;
    sine[1589]=662;
    sine[1590]=661;
    sine[1591]=660;
    sine[1592]=659;
    sine[1593]=658;
    sine[1594]=656;
    sine[1595]=655;
    sine[1596]=654;
    sine[1597]=653;
    sine[1598]=652;
    sine[1599]=650;
    sine[1600]=649;
    sine[1601]=648;
    sine[1602]=647;
    sine[1603]=645;
    sine[1604]=644;
    sine[1605]=643;
    sine[1606]=642;
    sine[1607]=641;
    sine[1608]=639;
    sine[1609]=638;
    sine[1610]=637;
    sine[1611]=636;
    sine[1612]=634;
    sine[1613]=633;
    sine[1614]=632;
    sine[1615]=631;
    sine[1616]=629;
    sine[1617]=628;
    sine[1618]=627;
    sine[1619]=626;
    sine[1620]=625;
    sine[1621]=623;
    sine[1622]=622;
    sine[1623]=621;
    sine[1624]=620;
    sine[1625]=618;
    sine[1626]=617;
    sine[1627]=616;
    sine[1628]=615;
    sine[1629]=613;
    sine[1630]=612;
    sine[1631]=611;
    sine[1632]=609;
    sine[1633]=608;
    sine[1634]=607;
    sine[1635]=606;
    sine[1636]=604;
    sine[1637]=603;
    sine[1638]=602;
    sine[1639]=601;
    sine[1640]=599;
    sine[1641]=598;
    sine[1642]=597;
    sine[1643]=596;
    sine[1644]=594;
    sine[1645]=593;
    sine[1646]=592;
    sine[1647]=590;
    sine[1648]=589;
    sine[1649]=588;
    sine[1650]=587;
    sine[1651]=585;
    sine[1652]=584;
    sine[1653]=583;
    sine[1654]=581;
    sine[1655]=580;
    sine[1656]=579;
    sine[1657]=578;
    sine[1658]=576;
    sine[1659]=575;
    sine[1660]=574;
    sine[1661]=572;
    sine[1662]=571;
    sine[1663]=570;
    sine[1664]=568;
    sine[1665]=567;
    sine[1666]=566;
    sine[1667]=564;
    sine[1668]=563;
    sine[1669]=562;
    sine[1670]=561;
    sine[1671]=559;
    sine[1672]=558;
    sine[1673]=557;
    sine[1674]=555;
    sine[1675]=554;
    sine[1676]=553;
    sine[1677]=551;
    sine[1678]=550;
    sine[1679]=549;
    sine[1680]=547;
    sine[1681]=546;
    sine[1682]=545;
    sine[1683]=543;
    sine[1684]=542;
    sine[1685]=541;
    sine[1686]=539;
    sine[1687]=538;
    sine[1688]=537;
    sine[1689]=535;
    sine[1690]=534;
    sine[1691]=533;
    sine[1692]=531;
    sine[1693]=530;
    sine[1694]=529;
    sine[1695]=527;
    sine[1696]=526;
    sine[1697]=525;
    sine[1698]=523;
    sine[1699]=522;
    sine[1700]=521;
    sine[1701]=519;
    sine[1702]=518;
    sine[1703]=516;
    sine[1704]=515;
    sine[1705]=514;
    sine[1706]=512;
    sine[1707]=511;
    sine[1708]=510;
    sine[1709]=508;
    sine[1710]=507;
    sine[1711]=506;
    sine[1712]=504;
    sine[1713]=503;
    sine[1714]=501;
    sine[1715]=500;
    sine[1716]=499;
    sine[1717]=497;
    sine[1718]=496;
    sine[1719]=495;
    sine[1720]=493;
    sine[1721]=492;
    sine[1722]=491;
    sine[1723]=489;
    sine[1724]=488;
    sine[1725]=486;
    sine[1726]=485;
    sine[1727]=484;
    sine[1728]=482;
    sine[1729]=481;
    sine[1730]=479;
    sine[1731]=478;
    sine[1732]=477;
    sine[1733]=475;
    sine[1734]=474;
    sine[1735]=472;
    sine[1736]=471;
    sine[1737]=470;
    sine[1738]=468;
    sine[1739]=467;
    sine[1740]=466;
    sine[1741]=464;
    sine[1742]=463;
    sine[1743]=461;
    sine[1744]=460;
    sine[1745]=458;
    sine[1746]=457;
    sine[1747]=456;
    sine[1748]=454;
    sine[1749]=453;
    sine[1750]=451;
    sine[1751]=450;
    sine[1752]=449;
    sine[1753]=447;
    sine[1754]=446;
    sine[1755]=444;
    sine[1756]=443;
    sine[1757]=442;
    sine[1758]=440;
    sine[1759]=439;
    sine[1760]=437;
    sine[1761]=436;
    sine[1762]=434;
    sine[1763]=433;
    sine[1764]=432;
    sine[1765]=430;
    sine[1766]=429;
    sine[1767]=427;
    sine[1768]=426;
    sine[1769]=424;
    sine[1770]=423;
    sine[1771]=422;
    sine[1772]=420;
    sine[1773]=419;
    sine[1774]=417;
    sine[1775]=416;
    sine[1776]=414;
    sine[1777]=413;
    sine[1778]=412;
    sine[1779]=410;
    sine[1780]=409;
    sine[1781]=407;
    sine[1782]=406;
    sine[1783]=404;
    sine[1784]=403;
    sine[1785]=402;
    sine[1786]=400;
    sine[1787]=399;
    sine[1788]=397;
    sine[1789]=396;
    sine[1790]=394;
    sine[1791]=393;
    sine[1792]=391;
    sine[1793]=390;
    sine[1794]=388;
    sine[1795]=387;
    sine[1796]=386;
    sine[1797]=384;
    sine[1798]=383;
    sine[1799]=381;
    sine[1800]=380;
    sine[1801]=378;
    sine[1802]=377;
    sine[1803]=375;
    sine[1804]=374;
    sine[1805]=372;
    sine[1806]=371;
    sine[1807]=369;
    sine[1808]=368;
    sine[1809]=367;
    sine[1810]=365;
    sine[1811]=364;
    sine[1812]=362;
    sine[1813]=361;
    sine[1814]=359;
    sine[1815]=358;
    sine[1816]=356;
    sine[1817]=355;
    sine[1818]=353;
    sine[1819]=352;
    sine[1820]=350;
    sine[1821]=349;
    sine[1822]=347;
    sine[1823]=346;
    sine[1824]=344;
    sine[1825]=343;
    sine[1826]=342;
    sine[1827]=340;
    sine[1828]=339;
    sine[1829]=337;
    sine[1830]=336;
    sine[1831]=334;
    sine[1832]=333;
    sine[1833]=331;
    sine[1834]=330;
    sine[1835]=328;
    sine[1836]=327;
    sine[1837]=325;
    sine[1838]=324;
    sine[1839]=322;
    sine[1840]=321;
    sine[1841]=319;
    sine[1842]=318;
    sine[1843]=316;
    sine[1844]=315;
    sine[1845]=313;
    sine[1846]=312;
    sine[1847]=310;
    sine[1848]=309;
    sine[1849]=307;
    sine[1850]=306;
    sine[1851]=304;
    sine[1852]=303;
    sine[1853]=301;
    sine[1854]=300;
    sine[1855]=298;
    sine[1856]=297;
    sine[1857]=295;
    sine[1858]=294;
    sine[1859]=292;
    sine[1860]=291;
    sine[1861]=289;
    sine[1862]=288;
    sine[1863]=286;
    sine[1864]=285;
    sine[1865]=283;
    sine[1866]=282;
    sine[1867]=280;
    sine[1868]=279;
    sine[1869]=277;
    sine[1870]=276;
    sine[1871]=274;
    sine[1872]=273;
    sine[1873]=271;
    sine[1874]=270;
    sine[1875]=268;
    sine[1876]=267;
    sine[1877]=265;
    sine[1878]=264;
    sine[1879]=262;
    sine[1880]=260;
    sine[1881]=259;
    sine[1882]=257;
    sine[1883]=256;
    sine[1884]=254;
    sine[1885]=253;
    sine[1886]=251;
    sine[1887]=250;
    sine[1888]=248;
    sine[1889]=247;
    sine[1890]=245;
    sine[1891]=244;
    sine[1892]=242;
    sine[1893]=241;
    sine[1894]=239;
    sine[1895]=238;
    sine[1896]=236;
    sine[1897]=235;
    sine[1898]=233;
    sine[1899]=232;
    sine[1900]=230;
    sine[1901]=228;
    sine[1902]=227;
    sine[1903]=225;
    sine[1904]=224;
    sine[1905]=222;
    sine[1906]=221;
    sine[1907]=219;
    sine[1908]=218;
    sine[1909]=216;
    sine[1910]=215;
    sine[1911]=213;
    sine[1912]=212;
    sine[1913]=210;
    sine[1914]=209;
    sine[1915]=207;
    sine[1916]=205;
    sine[1917]=204;
    sine[1918]=202;
    sine[1919]=201;
    sine[1920]=199;
    sine[1921]=198;
    sine[1922]=196;
    sine[1923]=195;
    sine[1924]=193;
    sine[1925]=192;
    sine[1926]=190;
    sine[1927]=188;
    sine[1928]=187;
    sine[1929]=185;
    sine[1930]=184;
    sine[1931]=182;
    sine[1932]=181;
    sine[1933]=179;
    sine[1934]=178;
    sine[1935]=176;
    sine[1936]=175;
    sine[1937]=173;
    sine[1938]=171;
    sine[1939]=170;
    sine[1940]=168;
    sine[1941]=167;
    sine[1942]=165;
    sine[1943]=164;
    sine[1944]=162;
    sine[1945]=161;
    sine[1946]=159;
    sine[1947]=158;
    sine[1948]=156;
    sine[1949]=154;
    sine[1950]=153;
    sine[1951]=151;
    sine[1952]=150;
    sine[1953]=148;
    sine[1954]=147;
    sine[1955]=145;
    sine[1956]=144;
    sine[1957]=142;
    sine[1958]=140;
    sine[1959]=139;
    sine[1960]=137;
    sine[1961]=136;
    sine[1962]=134;
    sine[1963]=133;
    sine[1964]=131;
    sine[1965]=130;
    sine[1966]=128;
    sine[1967]=126;
    sine[1968]=125;
    sine[1969]=123;
    sine[1970]=122;
    sine[1971]=120;
    sine[1972]=119;
    sine[1973]=117;
    sine[1974]=115;
    sine[1975]=114;
    sine[1976]=112;
    sine[1977]=111;
    sine[1978]=109;
    sine[1979]=108;
    sine[1980]=106;
    sine[1981]=105;
    sine[1982]=103;
    sine[1983]=101;
    sine[1984]=100;
    sine[1985]=98;
    sine[1986]=97;
    sine[1987]=95;
    sine[1988]=94;
    sine[1989]=92;
    sine[1990]=90;
    sine[1991]=89;
    sine[1992]=87;
    sine[1993]=86;
    sine[1994]=84;
    sine[1995]=83;
    sine[1996]=81;
    sine[1997]=80;
    sine[1998]=78;
    sine[1999]=76;
    sine[2000]=75;
    sine[2001]=73;
    sine[2002]=72;
    sine[2003]=70;
    sine[2004]=69;
    sine[2005]=67;
    sine[2006]=65;
    sine[2007]=64;
    sine[2008]=62;
    sine[2009]=61;
    sine[2010]=59;
    sine[2011]=58;
    sine[2012]=56;
    sine[2013]=54;
    sine[2014]=53;
    sine[2015]=51;
    sine[2016]=50;
    sine[2017]=48;
    sine[2018]=47;
    sine[2019]=45;
    sine[2020]=43;
    sine[2021]=42;
    sine[2022]=40;
    sine[2023]=39;
    sine[2024]=37;
    sine[2025]=36;
    sine[2026]=34;
    sine[2027]=32;
    sine[2028]=31;
    sine[2029]=29;
    sine[2030]=28;
    sine[2031]=26;
    sine[2032]=25;
    sine[2033]=23;
    sine[2034]=21;
    sine[2035]=20;
    sine[2036]=18;
    sine[2037]=17;
    sine[2038]=15;
    sine[2039]=14;
    sine[2040]=12;
    sine[2041]=10;
    sine[2042]=9;
    sine[2043]=7;
    sine[2044]=6;
    sine[2045]=4;
    sine[2046]=3;
    sine[2047]=1;
    sine[2048]=0;
    sine[2049]=-1;
    sine[2050]=-3;
    sine[2051]=-4;
    sine[2052]=-6;
    sine[2053]=-7;
    sine[2054]=-9;
    sine[2055]=-10;
    sine[2056]=-12;
    sine[2057]=-14;
    sine[2058]=-15;
    sine[2059]=-17;
    sine[2060]=-18;
    sine[2061]=-20;
    sine[2062]=-21;
    sine[2063]=-23;
    sine[2064]=-25;
    sine[2065]=-26;
    sine[2066]=-28;
    sine[2067]=-29;
    sine[2068]=-31;
    sine[2069]=-32;
    sine[2070]=-34;
    sine[2071]=-36;
    sine[2072]=-37;
    sine[2073]=-39;
    sine[2074]=-40;
    sine[2075]=-42;
    sine[2076]=-43;
    sine[2077]=-45;
    sine[2078]=-47;
    sine[2079]=-48;
    sine[2080]=-50;
    sine[2081]=-51;
    sine[2082]=-53;
    sine[2083]=-54;
    sine[2084]=-56;
    sine[2085]=-58;
    sine[2086]=-59;
    sine[2087]=-61;
    sine[2088]=-62;
    sine[2089]=-64;
    sine[2090]=-65;
    sine[2091]=-67;
    sine[2092]=-69;
    sine[2093]=-70;
    sine[2094]=-72;
    sine[2095]=-73;
    sine[2096]=-75;
    sine[2097]=-76;
    sine[2098]=-78;
    sine[2099]=-80;
    sine[2100]=-81;
    sine[2101]=-83;
    sine[2102]=-84;
    sine[2103]=-86;
    sine[2104]=-87;
    sine[2105]=-89;
    sine[2106]=-90;
    sine[2107]=-92;
    sine[2108]=-94;
    sine[2109]=-95;
    sine[2110]=-97;
    sine[2111]=-98;
    sine[2112]=-100;
    sine[2113]=-101;
    sine[2114]=-103;
    sine[2115]=-105;
    sine[2116]=-106;
    sine[2117]=-108;
    sine[2118]=-109;
    sine[2119]=-111;
    sine[2120]=-112;
    sine[2121]=-114;
    sine[2122]=-115;
    sine[2123]=-117;
    sine[2124]=-119;
    sine[2125]=-120;
    sine[2126]=-122;
    sine[2127]=-123;
    sine[2128]=-125;
    sine[2129]=-126;
    sine[2130]=-128;
    sine[2131]=-130;
    sine[2132]=-131;
    sine[2133]=-133;
    sine[2134]=-134;
    sine[2135]=-136;
    sine[2136]=-137;
    sine[2137]=-139;
    sine[2138]=-140;
    sine[2139]=-142;
    sine[2140]=-144;
    sine[2141]=-145;
    sine[2142]=-147;
    sine[2143]=-148;
    sine[2144]=-150;
    sine[2145]=-151;
    sine[2146]=-153;
    sine[2147]=-154;
    sine[2148]=-156;
    sine[2149]=-158;
    sine[2150]=-159;
    sine[2151]=-161;
    sine[2152]=-162;
    sine[2153]=-164;
    sine[2154]=-165;
    sine[2155]=-167;
    sine[2156]=-168;
    sine[2157]=-170;
    sine[2158]=-171;
    sine[2159]=-173;
    sine[2160]=-175;
    sine[2161]=-176;
    sine[2162]=-178;
    sine[2163]=-179;
    sine[2164]=-181;
    sine[2165]=-182;
    sine[2166]=-184;
    sine[2167]=-185;
    sine[2168]=-187;
    sine[2169]=-188;
    sine[2170]=-190;
    sine[2171]=-192;
    sine[2172]=-193;
    sine[2173]=-195;
    sine[2174]=-196;
    sine[2175]=-198;
    sine[2176]=-199;
    sine[2177]=-201;
    sine[2178]=-202;
    sine[2179]=-204;
    sine[2180]=-205;
    sine[2181]=-207;
    sine[2182]=-209;
    sine[2183]=-210;
    sine[2184]=-212;
    sine[2185]=-213;
    sine[2186]=-215;
    sine[2187]=-216;
    sine[2188]=-218;
    sine[2189]=-219;
    sine[2190]=-221;
    sine[2191]=-222;
    sine[2192]=-224;
    sine[2193]=-225;
    sine[2194]=-227;
    sine[2195]=-228;
    sine[2196]=-230;
    sine[2197]=-232;
    sine[2198]=-233;
    sine[2199]=-235;
    sine[2200]=-236;
    sine[2201]=-238;
    sine[2202]=-239;
    sine[2203]=-241;
    sine[2204]=-242;
    sine[2205]=-244;
    sine[2206]=-245;
    sine[2207]=-247;
    sine[2208]=-248;
    sine[2209]=-250;
    sine[2210]=-251;
    sine[2211]=-253;
    sine[2212]=-254;
    sine[2213]=-256;
    sine[2214]=-257;
    sine[2215]=-259;
    sine[2216]=-260;
    sine[2217]=-262;
    sine[2218]=-264;
    sine[2219]=-265;
    sine[2220]=-267;
    sine[2221]=-268;
    sine[2222]=-270;
    sine[2223]=-271;
    sine[2224]=-273;
    sine[2225]=-274;
    sine[2226]=-276;
    sine[2227]=-277;
    sine[2228]=-279;
    sine[2229]=-280;
    sine[2230]=-282;
    sine[2231]=-283;
    sine[2232]=-285;
    sine[2233]=-286;
    sine[2234]=-288;
    sine[2235]=-289;
    sine[2236]=-291;
    sine[2237]=-292;
    sine[2238]=-294;
    sine[2239]=-295;
    sine[2240]=-297;
    sine[2241]=-298;
    sine[2242]=-300;
    sine[2243]=-301;
    sine[2244]=-303;
    sine[2245]=-304;
    sine[2246]=-306;
    sine[2247]=-307;
    sine[2248]=-309;
    sine[2249]=-310;
    sine[2250]=-312;
    sine[2251]=-313;
    sine[2252]=-315;
    sine[2253]=-316;
    sine[2254]=-318;
    sine[2255]=-319;
    sine[2256]=-321;
    sine[2257]=-322;
    sine[2258]=-324;
    sine[2259]=-325;
    sine[2260]=-327;
    sine[2261]=-328;
    sine[2262]=-330;
    sine[2263]=-331;
    sine[2264]=-333;
    sine[2265]=-334;
    sine[2266]=-336;
    sine[2267]=-337;
    sine[2268]=-339;
    sine[2269]=-340;
    sine[2270]=-342;
    sine[2271]=-343;
    sine[2272]=-344;
    sine[2273]=-346;
    sine[2274]=-347;
    sine[2275]=-349;
    sine[2276]=-350;
    sine[2277]=-352;
    sine[2278]=-353;
    sine[2279]=-355;
    sine[2280]=-356;
    sine[2281]=-358;
    sine[2282]=-359;
    sine[2283]=-361;
    sine[2284]=-362;
    sine[2285]=-364;
    sine[2286]=-365;
    sine[2287]=-367;
    sine[2288]=-368;
    sine[2289]=-369;
    sine[2290]=-371;
    sine[2291]=-372;
    sine[2292]=-374;
    sine[2293]=-375;
    sine[2294]=-377;
    sine[2295]=-378;
    sine[2296]=-380;
    sine[2297]=-381;
    sine[2298]=-383;
    sine[2299]=-384;
    sine[2300]=-386;
    sine[2301]=-387;
    sine[2302]=-388;
    sine[2303]=-390;
    sine[2304]=-391;
    sine[2305]=-393;
    sine[2306]=-394;
    sine[2307]=-396;
    sine[2308]=-397;
    sine[2309]=-399;
    sine[2310]=-400;
    sine[2311]=-402;
    sine[2312]=-403;
    sine[2313]=-404;
    sine[2314]=-406;
    sine[2315]=-407;
    sine[2316]=-409;
    sine[2317]=-410;
    sine[2318]=-412;
    sine[2319]=-413;
    sine[2320]=-414;
    sine[2321]=-416;
    sine[2322]=-417;
    sine[2323]=-419;
    sine[2324]=-420;
    sine[2325]=-422;
    sine[2326]=-423;
    sine[2327]=-424;
    sine[2328]=-426;
    sine[2329]=-427;
    sine[2330]=-429;
    sine[2331]=-430;
    sine[2332]=-432;
    sine[2333]=-433;
    sine[2334]=-434;
    sine[2335]=-436;
    sine[2336]=-437;
    sine[2337]=-439;
    sine[2338]=-440;
    sine[2339]=-442;
    sine[2340]=-443;
    sine[2341]=-444;
    sine[2342]=-446;
    sine[2343]=-447;
    sine[2344]=-449;
    sine[2345]=-450;
    sine[2346]=-451;
    sine[2347]=-453;
    sine[2348]=-454;
    sine[2349]=-456;
    sine[2350]=-457;
    sine[2351]=-458;
    sine[2352]=-460;
    sine[2353]=-461;
    sine[2354]=-463;
    sine[2355]=-464;
    sine[2356]=-466;
    sine[2357]=-467;
    sine[2358]=-468;
    sine[2359]=-470;
    sine[2360]=-471;
    sine[2361]=-472;
    sine[2362]=-474;
    sine[2363]=-475;
    sine[2364]=-477;
    sine[2365]=-478;
    sine[2366]=-479;
    sine[2367]=-481;
    sine[2368]=-482;
    sine[2369]=-484;
    sine[2370]=-485;
    sine[2371]=-486;
    sine[2372]=-488;
    sine[2373]=-489;
    sine[2374]=-491;
    sine[2375]=-492;
    sine[2376]=-493;
    sine[2377]=-495;
    sine[2378]=-496;
    sine[2379]=-497;
    sine[2380]=-499;
    sine[2381]=-500;
    sine[2382]=-501;
    sine[2383]=-503;
    sine[2384]=-504;
    sine[2385]=-506;
    sine[2386]=-507;
    sine[2387]=-508;
    sine[2388]=-510;
    sine[2389]=-511;
    sine[2390]=-512;
    sine[2391]=-514;
    sine[2392]=-515;
    sine[2393]=-516;
    sine[2394]=-518;
    sine[2395]=-519;
    sine[2396]=-521;
    sine[2397]=-522;
    sine[2398]=-523;
    sine[2399]=-525;
    sine[2400]=-526;
    sine[2401]=-527;
    sine[2402]=-529;
    sine[2403]=-530;
    sine[2404]=-531;
    sine[2405]=-533;
    sine[2406]=-534;
    sine[2407]=-535;
    sine[2408]=-537;
    sine[2409]=-538;
    sine[2410]=-539;
    sine[2411]=-541;
    sine[2412]=-542;
    sine[2413]=-543;
    sine[2414]=-545;
    sine[2415]=-546;
    sine[2416]=-547;
    sine[2417]=-549;
    sine[2418]=-550;
    sine[2419]=-551;
    sine[2420]=-553;
    sine[2421]=-554;
    sine[2422]=-555;
    sine[2423]=-557;
    sine[2424]=-558;
    sine[2425]=-559;
    sine[2426]=-561;
    sine[2427]=-562;
    sine[2428]=-563;
    sine[2429]=-564;
    sine[2430]=-566;
    sine[2431]=-567;
    sine[2432]=-568;
    sine[2433]=-570;
    sine[2434]=-571;
    sine[2435]=-572;
    sine[2436]=-574;
    sine[2437]=-575;
    sine[2438]=-576;
    sine[2439]=-578;
    sine[2440]=-579;
    sine[2441]=-580;
    sine[2442]=-581;
    sine[2443]=-583;
    sine[2444]=-584;
    sine[2445]=-585;
    sine[2446]=-587;
    sine[2447]=-588;
    sine[2448]=-589;
    sine[2449]=-590;
    sine[2450]=-592;
    sine[2451]=-593;
    sine[2452]=-594;
    sine[2453]=-596;
    sine[2454]=-597;
    sine[2455]=-598;
    sine[2456]=-599;
    sine[2457]=-601;
    sine[2458]=-602;
    sine[2459]=-603;
    sine[2460]=-604;
    sine[2461]=-606;
    sine[2462]=-607;
    sine[2463]=-608;
    sine[2464]=-609;
    sine[2465]=-611;
    sine[2466]=-612;
    sine[2467]=-613;
    sine[2468]=-615;
    sine[2469]=-616;
    sine[2470]=-617;
    sine[2471]=-618;
    sine[2472]=-620;
    sine[2473]=-621;
    sine[2474]=-622;
    sine[2475]=-623;
    sine[2476]=-625;
    sine[2477]=-626;
    sine[2478]=-627;
    sine[2479]=-628;
    sine[2480]=-629;
    sine[2481]=-631;
    sine[2482]=-632;
    sine[2483]=-633;
    sine[2484]=-634;
    sine[2485]=-636;
    sine[2486]=-637;
    sine[2487]=-638;
    sine[2488]=-639;
    sine[2489]=-641;
    sine[2490]=-642;
    sine[2491]=-643;
    sine[2492]=-644;
    sine[2493]=-645;
    sine[2494]=-647;
    sine[2495]=-648;
    sine[2496]=-649;
    sine[2497]=-650;
    sine[2498]=-652;
    sine[2499]=-653;
    sine[2500]=-654;
    sine[2501]=-655;
    sine[2502]=-656;
    sine[2503]=-658;
    sine[2504]=-659;
    sine[2505]=-660;
    sine[2506]=-661;
    sine[2507]=-662;
    sine[2508]=-664;
    sine[2509]=-665;
    sine[2510]=-666;
    sine[2511]=-667;
    sine[2512]=-668;
    sine[2513]=-670;
    sine[2514]=-671;
    sine[2515]=-672;
    sine[2516]=-673;
    sine[2517]=-674;
    sine[2518]=-675;
    sine[2519]=-677;
    sine[2520]=-678;
    sine[2521]=-679;
    sine[2522]=-680;
    sine[2523]=-681;
    sine[2524]=-683;
    sine[2525]=-684;
    sine[2526]=-685;
    sine[2527]=-686;
    sine[2528]=-687;
    sine[2529]=-688;
    sine[2530]=-690;
    sine[2531]=-691;
    sine[2532]=-692;
    sine[2533]=-693;
    sine[2534]=-694;
    sine[2535]=-695;
    sine[2536]=-696;
    sine[2537]=-698;
    sine[2538]=-699;
    sine[2539]=-700;
    sine[2540]=-701;
    sine[2541]=-702;
    sine[2542]=-703;
    sine[2543]=-704;
    sine[2544]=-706;
    sine[2545]=-707;
    sine[2546]=-708;
    sine[2547]=-709;
    sine[2548]=-710;
    sine[2549]=-711;
    sine[2550]=-712;
    sine[2551]=-714;
    sine[2552]=-715;
    sine[2553]=-716;
    sine[2554]=-717;
    sine[2555]=-718;
    sine[2556]=-719;
    sine[2557]=-720;
    sine[2558]=-721;
    sine[2559]=-722;
    sine[2560]=-724;
    sine[2561]=-725;
    sine[2562]=-726;
    sine[2563]=-727;
    sine[2564]=-728;
    sine[2565]=-729;
    sine[2566]=-730;
    sine[2567]=-731;
    sine[2568]=-732;
    sine[2569]=-734;
    sine[2570]=-735;
    sine[2571]=-736;
    sine[2572]=-737;
    sine[2573]=-738;
    sine[2574]=-739;
    sine[2575]=-740;
    sine[2576]=-741;
    sine[2577]=-742;
    sine[2578]=-743;
    sine[2579]=-744;
    sine[2580]=-745;
    sine[2581]=-747;
    sine[2582]=-748;
    sine[2583]=-749;
    sine[2584]=-750;
    sine[2585]=-751;
    sine[2586]=-752;
    sine[2587]=-753;
    sine[2588]=-754;
    sine[2589]=-755;
    sine[2590]=-756;
    sine[2591]=-757;
    sine[2592]=-758;
    sine[2593]=-759;
    sine[2594]=-760;
    sine[2595]=-761;
    sine[2596]=-762;
    sine[2597]=-763;
    sine[2598]=-765;
    sine[2599]=-766;
    sine[2600]=-767;
    sine[2601]=-768;
    sine[2602]=-769;
    sine[2603]=-770;
    sine[2604]=-771;
    sine[2605]=-772;
    sine[2606]=-773;
    sine[2607]=-774;
    sine[2608]=-775;
    sine[2609]=-776;
    sine[2610]=-777;
    sine[2611]=-778;
    sine[2612]=-779;
    sine[2613]=-780;
    sine[2614]=-781;
    sine[2615]=-782;
    sine[2616]=-783;
    sine[2617]=-784;
    sine[2618]=-785;
    sine[2619]=-786;
    sine[2620]=-787;
    sine[2621]=-788;
    sine[2622]=-789;
    sine[2623]=-790;
    sine[2624]=-791;
    sine[2625]=-792;
    sine[2626]=-793;
    sine[2627]=-794;
    sine[2628]=-795;
    sine[2629]=-796;
    sine[2630]=-797;
    sine[2631]=-798;
    sine[2632]=-799;
    sine[2633]=-800;
    sine[2634]=-801;
    sine[2635]=-802;
    sine[2636]=-803;
    sine[2637]=-804;
    sine[2638]=-805;
    sine[2639]=-806;
    sine[2640]=-807;
    sine[2641]=-808;
    sine[2642]=-809;
    sine[2643]=-810;
    sine[2644]=-811;
    sine[2645]=-812;
    sine[2646]=-813;
    sine[2647]=-813;
    sine[2648]=-814;
    sine[2649]=-815;
    sine[2650]=-816;
    sine[2651]=-817;
    sine[2652]=-818;
    sine[2653]=-819;
    sine[2654]=-820;
    sine[2655]=-821;
    sine[2656]=-822;
    sine[2657]=-823;
    sine[2658]=-824;
    sine[2659]=-825;
    sine[2660]=-826;
    sine[2661]=-827;
    sine[2662]=-828;
    sine[2663]=-828;
    sine[2664]=-829;
    sine[2665]=-830;
    sine[2666]=-831;
    sine[2667]=-832;
    sine[2668]=-833;
    sine[2669]=-834;
    sine[2670]=-835;
    sine[2671]=-836;
    sine[2672]=-837;
    sine[2673]=-838;
    sine[2674]=-839;
    sine[2675]=-839;
    sine[2676]=-840;
    sine[2677]=-841;
    sine[2678]=-842;
    sine[2679]=-843;
    sine[2680]=-844;
    sine[2681]=-845;
    sine[2682]=-846;
    sine[2683]=-847;
    sine[2684]=-847;
    sine[2685]=-848;
    sine[2686]=-849;
    sine[2687]=-850;
    sine[2688]=-851;
    sine[2689]=-852;
    sine[2690]=-853;
    sine[2691]=-854;
    sine[2692]=-854;
    sine[2693]=-855;
    sine[2694]=-856;
    sine[2695]=-857;
    sine[2696]=-858;
    sine[2697]=-859;
    sine[2698]=-860;
    sine[2699]=-860;
    sine[2700]=-861;
    sine[2701]=-862;
    sine[2702]=-863;
    sine[2703]=-864;
    sine[2704]=-865;
    sine[2705]=-865;
    sine[2706]=-866;
    sine[2707]=-867;
    sine[2708]=-868;
    sine[2709]=-869;
    sine[2710]=-870;
    sine[2711]=-870;
    sine[2712]=-871;
    sine[2713]=-872;
    sine[2714]=-873;
    sine[2715]=-874;
    sine[2716]=-875;
    sine[2717]=-875;
    sine[2718]=-876;
    sine[2719]=-877;
    sine[2720]=-878;
    sine[2721]=-879;
    sine[2722]=-879;
    sine[2723]=-880;
    sine[2724]=-881;
    sine[2725]=-882;
    sine[2726]=-883;
    sine[2727]=-883;
    sine[2728]=-884;
    sine[2729]=-885;
    sine[2730]=-886;
    sine[2731]=-887;
    sine[2732]=-887;
    sine[2733]=-888;
    sine[2734]=-889;
    sine[2735]=-890;
    sine[2736]=-890;
    sine[2737]=-891;
    sine[2738]=-892;
    sine[2739]=-893;
    sine[2740]=-894;
    sine[2741]=-894;
    sine[2742]=-895;
    sine[2743]=-896;
    sine[2744]=-897;
    sine[2745]=-897;
    sine[2746]=-898;
    sine[2747]=-899;
    sine[2748]=-900;
    sine[2749]=-900;
    sine[2750]=-901;
    sine[2751]=-902;
    sine[2752]=-903;
    sine[2753]=-903;
    sine[2754]=-904;
    sine[2755]=-905;
    sine[2756]=-906;
    sine[2757]=-906;
    sine[2758]=-907;
    sine[2759]=-908;
    sine[2760]=-908;
    sine[2761]=-909;
    sine[2762]=-910;
    sine[2763]=-911;
    sine[2764]=-911;
    sine[2765]=-912;
    sine[2766]=-913;
    sine[2767]=-913;
    sine[2768]=-914;
    sine[2769]=-915;
    sine[2770]=-916;
    sine[2771]=-916;
    sine[2772]=-917;
    sine[2773]=-918;
    sine[2774]=-918;
    sine[2775]=-919;
    sine[2776]=-920;
    sine[2777]=-920;
    sine[2778]=-921;
    sine[2779]=-922;
    sine[2780]=-922;
    sine[2781]=-923;
    sine[2782]=-924;
    sine[2783]=-925;
    sine[2784]=-925;
    sine[2785]=-926;
    sine[2786]=-927;
    sine[2787]=-927;
    sine[2788]=-928;
    sine[2789]=-929;
    sine[2790]=-929;
    sine[2791]=-930;
    sine[2792]=-930;
    sine[2793]=-931;
    sine[2794]=-932;
    sine[2795]=-932;
    sine[2796]=-933;
    sine[2797]=-934;
    sine[2798]=-934;
    sine[2799]=-935;
    sine[2800]=-936;
    sine[2801]=-936;
    sine[2802]=-937;
    sine[2803]=-938;
    sine[2804]=-938;
    sine[2805]=-939;
    sine[2806]=-939;
    sine[2807]=-940;
    sine[2808]=-941;
    sine[2809]=-941;
    sine[2810]=-942;
    sine[2811]=-943;
    sine[2812]=-943;
    sine[2813]=-944;
    sine[2814]=-944;
    sine[2815]=-945;
    sine[2816]=-946;
    sine[2817]=-946;
    sine[2818]=-947;
    sine[2819]=-947;
    sine[2820]=-948;
    sine[2821]=-949;
    sine[2822]=-949;
    sine[2823]=-950;
    sine[2824]=-950;
    sine[2825]=-951;
    sine[2826]=-951;
    sine[2827]=-952;
    sine[2828]=-953;
    sine[2829]=-953;
    sine[2830]=-954;
    sine[2831]=-954;
    sine[2832]=-955;
    sine[2833]=-955;
    sine[2834]=-956;
    sine[2835]=-957;
    sine[2836]=-957;
    sine[2837]=-958;
    sine[2838]=-958;
    sine[2839]=-959;
    sine[2840]=-959;
    sine[2841]=-960;
    sine[2842]=-960;
    sine[2843]=-961;
    sine[2844]=-962;
    sine[2845]=-962;
    sine[2846]=-963;
    sine[2847]=-963;
    sine[2848]=-964;
    sine[2849]=-964;
    sine[2850]=-965;
    sine[2851]=-965;
    sine[2852]=-966;
    sine[2853]=-966;
    sine[2854]=-967;
    sine[2855]=-967;
    sine[2856]=-968;
    sine[2857]=-968;
    sine[2858]=-969;
    sine[2859]=-969;
    sine[2860]=-970;
    sine[2861]=-970;
    sine[2862]=-971;
    sine[2863]=-971;
    sine[2864]=-972;
    sine[2865]=-972;
    sine[2866]=-973;
    sine[2867]=-973;
    sine[2868]=-974;
    sine[2869]=-974;
    sine[2870]=-975;
    sine[2871]=-975;
    sine[2872]=-976;
    sine[2873]=-976;
    sine[2874]=-977;
    sine[2875]=-977;
    sine[2876]=-978;
    sine[2877]=-978;
    sine[2878]=-978;
    sine[2879]=-979;
    sine[2880]=-979;
    sine[2881]=-980;
    sine[2882]=-980;
    sine[2883]=-981;
    sine[2884]=-981;
    sine[2885]=-982;
    sine[2886]=-982;
    sine[2887]=-983;
    sine[2888]=-983;
    sine[2889]=-983;
    sine[2890]=-984;
    sine[2891]=-984;
    sine[2892]=-985;
    sine[2893]=-985;
    sine[2894]=-986;
    sine[2895]=-986;
    sine[2896]=-986;
    sine[2897]=-987;
    sine[2898]=-987;
    sine[2899]=-988;
    sine[2900]=-988;
    sine[2901]=-988;
    sine[2902]=-989;
    sine[2903]=-989;
    sine[2904]=-990;
    sine[2905]=-990;
    sine[2906]=-990;
    sine[2907]=-991;
    sine[2908]=-991;
    sine[2909]=-992;
    sine[2910]=-992;
    sine[2911]=-992;
    sine[2912]=-993;
    sine[2913]=-993;
    sine[2914]=-994;
    sine[2915]=-994;
    sine[2916]=-994;
    sine[2917]=-995;
    sine[2918]=-995;
    sine[2919]=-995;
    sine[2920]=-996;
    sine[2921]=-996;
    sine[2922]=-997;
    sine[2923]=-997;
    sine[2924]=-997;
    sine[2925]=-998;
    sine[2926]=-998;
    sine[2927]=-998;
    sine[2928]=-999;
    sine[2929]=-999;
    sine[2930]=-999;
    sine[2931]=-1000;
    sine[2932]=-1000;
    sine[2933]=-1000;
    sine[2934]=-1001;
    sine[2935]=-1001;
    sine[2936]=-1001;
    sine[2937]=-1002;
    sine[2938]=-1002;
    sine[2939]=-1002;
    sine[2940]=-1003;
    sine[2941]=-1003;
    sine[2942]=-1003;
    sine[2943]=-1004;
    sine[2944]=-1004;
    sine[2945]=-1004;
    sine[2946]=-1004;
    sine[2947]=-1005;
    sine[2948]=-1005;
    sine[2949]=-1005;
    sine[2950]=-1006;
    sine[2951]=-1006;
    sine[2952]=-1006;
    sine[2953]=-1006;
    sine[2954]=-1007;
    sine[2955]=-1007;
    sine[2956]=-1007;
    sine[2957]=-1008;
    sine[2958]=-1008;
    sine[2959]=-1008;
    sine[2960]=-1008;
    sine[2961]=-1009;
    sine[2962]=-1009;
    sine[2963]=-1009;
    sine[2964]=-1009;
    sine[2965]=-1010;
    sine[2966]=-1010;
    sine[2967]=-1010;
    sine[2968]=-1010;
    sine[2969]=-1011;
    sine[2970]=-1011;
    sine[2971]=-1011;
    sine[2972]=-1011;
    sine[2973]=-1012;
    sine[2974]=-1012;
    sine[2975]=-1012;
    sine[2976]=-1012;
    sine[2977]=-1013;
    sine[2978]=-1013;
    sine[2979]=-1013;
    sine[2980]=-1013;
    sine[2981]=-1014;
    sine[2982]=-1014;
    sine[2983]=-1014;
    sine[2984]=-1014;
    sine[2985]=-1014;
    sine[2986]=-1015;
    sine[2987]=-1015;
    sine[2988]=-1015;
    sine[2989]=-1015;
    sine[2990]=-1015;
    sine[2991]=-1016;
    sine[2992]=-1016;
    sine[2993]=-1016;
    sine[2994]=-1016;
    sine[2995]=-1016;
    sine[2996]=-1017;
    sine[2997]=-1017;
    sine[2998]=-1017;
    sine[2999]=-1017;
    sine[3000]=-1017;
    sine[3001]=-1017;
    sine[3002]=-1018;
    sine[3003]=-1018;
    sine[3004]=-1018;
    sine[3005]=-1018;
    sine[3006]=-1018;
    sine[3007]=-1018;
    sine[3008]=-1019;
    sine[3009]=-1019;
    sine[3010]=-1019;
    sine[3011]=-1019;
    sine[3012]=-1019;
    sine[3013]=-1019;
    sine[3014]=-1019;
    sine[3015]=-1020;
    sine[3016]=-1020;
    sine[3017]=-1020;
    sine[3018]=-1020;
    sine[3019]=-1020;
    sine[3020]=-1020;
    sine[3021]=-1020;
    sine[3022]=-1020;
    sine[3023]=-1021;
    sine[3024]=-1021;
    sine[3025]=-1021;
    sine[3026]=-1021;
    sine[3027]=-1021;
    sine[3028]=-1021;
    sine[3029]=-1021;
    sine[3030]=-1021;
    sine[3031]=-1021;
    sine[3032]=-1022;
    sine[3033]=-1022;
    sine[3034]=-1022;
    sine[3035]=-1022;
    sine[3036]=-1022;
    sine[3037]=-1022;
    sine[3038]=-1022;
    sine[3039]=-1022;
    sine[3040]=-1022;
    sine[3041]=-1022;
    sine[3042]=-1022;
    sine[3043]=-1022;
    sine[3044]=-1023;
    sine[3045]=-1023;
    sine[3046]=-1023;
    sine[3047]=-1023;
    sine[3048]=-1023;
    sine[3049]=-1023;
    sine[3050]=-1023;
    sine[3051]=-1023;
    sine[3052]=-1023;
    sine[3053]=-1023;
    sine[3054]=-1023;
    sine[3055]=-1023;
    sine[3056]=-1023;
    sine[3057]=-1023;
    sine[3058]=-1023;
    sine[3059]=-1023;
    sine[3060]=-1023;
    sine[3061]=-1023;
    sine[3062]=-1023;
    sine[3063]=-1023;
    sine[3064]=-1023;
    sine[3065]=-1023;
    sine[3066]=-1023;
    sine[3067]=-1023;
    sine[3068]=-1023;
    sine[3069]=-1023;
    sine[3070]=-1023;
    sine[3071]=-1023;
    sine[3072]=-1024;
    sine[3073]=-1023;
    sine[3074]=-1023;
    sine[3075]=-1023;
    sine[3076]=-1023;
    sine[3077]=-1023;
    sine[3078]=-1023;
    sine[3079]=-1023;
    sine[3080]=-1023;
    sine[3081]=-1023;
    sine[3082]=-1023;
    sine[3083]=-1023;
    sine[3084]=-1023;
    sine[3085]=-1023;
    sine[3086]=-1023;
    sine[3087]=-1023;
    sine[3088]=-1023;
    sine[3089]=-1023;
    sine[3090]=-1023;
    sine[3091]=-1023;
    sine[3092]=-1023;
    sine[3093]=-1023;
    sine[3094]=-1023;
    sine[3095]=-1023;
    sine[3096]=-1023;
    sine[3097]=-1023;
    sine[3098]=-1023;
    sine[3099]=-1023;
    sine[3100]=-1023;
    sine[3101]=-1022;
    sine[3102]=-1022;
    sine[3103]=-1022;
    sine[3104]=-1022;
    sine[3105]=-1022;
    sine[3106]=-1022;
    sine[3107]=-1022;
    sine[3108]=-1022;
    sine[3109]=-1022;
    sine[3110]=-1022;
    sine[3111]=-1022;
    sine[3112]=-1022;
    sine[3113]=-1021;
    sine[3114]=-1021;
    sine[3115]=-1021;
    sine[3116]=-1021;
    sine[3117]=-1021;
    sine[3118]=-1021;
    sine[3119]=-1021;
    sine[3120]=-1021;
    sine[3121]=-1021;
    sine[3122]=-1020;
    sine[3123]=-1020;
    sine[3124]=-1020;
    sine[3125]=-1020;
    sine[3126]=-1020;
    sine[3127]=-1020;
    sine[3128]=-1020;
    sine[3129]=-1020;
    sine[3130]=-1019;
    sine[3131]=-1019;
    sine[3132]=-1019;
    sine[3133]=-1019;
    sine[3134]=-1019;
    sine[3135]=-1019;
    sine[3136]=-1019;
    sine[3137]=-1018;
    sine[3138]=-1018;
    sine[3139]=-1018;
    sine[3140]=-1018;
    sine[3141]=-1018;
    sine[3142]=-1018;
    sine[3143]=-1017;
    sine[3144]=-1017;
    sine[3145]=-1017;
    sine[3146]=-1017;
    sine[3147]=-1017;
    sine[3148]=-1017;
    sine[3149]=-1016;
    sine[3150]=-1016;
    sine[3151]=-1016;
    sine[3152]=-1016;
    sine[3153]=-1016;
    sine[3154]=-1015;
    sine[3155]=-1015;
    sine[3156]=-1015;
    sine[3157]=-1015;
    sine[3158]=-1015;
    sine[3159]=-1014;
    sine[3160]=-1014;
    sine[3161]=-1014;
    sine[3162]=-1014;
    sine[3163]=-1014;
    sine[3164]=-1013;
    sine[3165]=-1013;
    sine[3166]=-1013;
    sine[3167]=-1013;
    sine[3168]=-1012;
    sine[3169]=-1012;
    sine[3170]=-1012;
    sine[3171]=-1012;
    sine[3172]=-1011;
    sine[3173]=-1011;
    sine[3174]=-1011;
    sine[3175]=-1011;
    sine[3176]=-1010;
    sine[3177]=-1010;
    sine[3178]=-1010;
    sine[3179]=-1010;
    sine[3180]=-1009;
    sine[3181]=-1009;
    sine[3182]=-1009;
    sine[3183]=-1009;
    sine[3184]=-1008;
    sine[3185]=-1008;
    sine[3186]=-1008;
    sine[3187]=-1008;
    sine[3188]=-1007;
    sine[3189]=-1007;
    sine[3190]=-1007;
    sine[3191]=-1006;
    sine[3192]=-1006;
    sine[3193]=-1006;
    sine[3194]=-1006;
    sine[3195]=-1005;
    sine[3196]=-1005;
    sine[3197]=-1005;
    sine[3198]=-1004;
    sine[3199]=-1004;
    sine[3200]=-1004;
    sine[3201]=-1004;
    sine[3202]=-1003;
    sine[3203]=-1003;
    sine[3204]=-1003;
    sine[3205]=-1002;
    sine[3206]=-1002;
    sine[3207]=-1002;
    sine[3208]=-1001;
    sine[3209]=-1001;
    sine[3210]=-1001;
    sine[3211]=-1000;
    sine[3212]=-1000;
    sine[3213]=-1000;
    sine[3214]=-999;
    sine[3215]=-999;
    sine[3216]=-999;
    sine[3217]=-998;
    sine[3218]=-998;
    sine[3219]=-998;
    sine[3220]=-997;
    sine[3221]=-997;
    sine[3222]=-997;
    sine[3223]=-996;
    sine[3224]=-996;
    sine[3225]=-995;
    sine[3226]=-995;
    sine[3227]=-995;
    sine[3228]=-994;
    sine[3229]=-994;
    sine[3230]=-994;
    sine[3231]=-993;
    sine[3232]=-993;
    sine[3233]=-992;
    sine[3234]=-992;
    sine[3235]=-992;
    sine[3236]=-991;
    sine[3237]=-991;
    sine[3238]=-990;
    sine[3239]=-990;
    sine[3240]=-990;
    sine[3241]=-989;
    sine[3242]=-989;
    sine[3243]=-988;
    sine[3244]=-988;
    sine[3245]=-988;
    sine[3246]=-987;
    sine[3247]=-987;
    sine[3248]=-986;
    sine[3249]=-986;
    sine[3250]=-986;
    sine[3251]=-985;
    sine[3252]=-985;
    sine[3253]=-984;
    sine[3254]=-984;
    sine[3255]=-983;
    sine[3256]=-983;
    sine[3257]=-983;
    sine[3258]=-982;
    sine[3259]=-982;
    sine[3260]=-981;
    sine[3261]=-981;
    sine[3262]=-980;
    sine[3263]=-980;
    sine[3264]=-979;
    sine[3265]=-979;
    sine[3266]=-978;
    sine[3267]=-978;
    sine[3268]=-978;
    sine[3269]=-977;
    sine[3270]=-977;
    sine[3271]=-976;
    sine[3272]=-976;
    sine[3273]=-975;
    sine[3274]=-975;
    sine[3275]=-974;
    sine[3276]=-974;
    sine[3277]=-973;
    sine[3278]=-973;
    sine[3279]=-972;
    sine[3280]=-972;
    sine[3281]=-971;
    sine[3282]=-971;
    sine[3283]=-970;
    sine[3284]=-970;
    sine[3285]=-969;
    sine[3286]=-969;
    sine[3287]=-968;
    sine[3288]=-968;
    sine[3289]=-967;
    sine[3290]=-967;
    sine[3291]=-966;
    sine[3292]=-966;
    sine[3293]=-965;
    sine[3294]=-965;
    sine[3295]=-964;
    sine[3296]=-964;
    sine[3297]=-963;
    sine[3298]=-963;
    sine[3299]=-962;
    sine[3300]=-962;
    sine[3301]=-961;
    sine[3302]=-960;
    sine[3303]=-960;
    sine[3304]=-959;
    sine[3305]=-959;
    sine[3306]=-958;
    sine[3307]=-958;
    sine[3308]=-957;
    sine[3309]=-957;
    sine[3310]=-956;
    sine[3311]=-955;
    sine[3312]=-955;
    sine[3313]=-954;
    sine[3314]=-954;
    sine[3315]=-953;
    sine[3316]=-953;
    sine[3317]=-952;
    sine[3318]=-951;
    sine[3319]=-951;
    sine[3320]=-950;
    sine[3321]=-950;
    sine[3322]=-949;
    sine[3323]=-949;
    sine[3324]=-948;
    sine[3325]=-947;
    sine[3326]=-947;
    sine[3327]=-946;
    sine[3328]=-946;
    sine[3329]=-945;
    sine[3330]=-944;
    sine[3331]=-944;
    sine[3332]=-943;
    sine[3333]=-943;
    sine[3334]=-942;
    sine[3335]=-941;
    sine[3336]=-941;
    sine[3337]=-940;
    sine[3338]=-939;
    sine[3339]=-939;
    sine[3340]=-938;
    sine[3341]=-938;
    sine[3342]=-937;
    sine[3343]=-936;
    sine[3344]=-936;
    sine[3345]=-935;
    sine[3346]=-934;
    sine[3347]=-934;
    sine[3348]=-933;
    sine[3349]=-932;
    sine[3350]=-932;
    sine[3351]=-931;
    sine[3352]=-930;
    sine[3353]=-930;
    sine[3354]=-929;
    sine[3355]=-929;
    sine[3356]=-928;
    sine[3357]=-927;
    sine[3358]=-927;
    sine[3359]=-926;
    sine[3360]=-925;
    sine[3361]=-925;
    sine[3362]=-924;
    sine[3363]=-923;
    sine[3364]=-922;
    sine[3365]=-922;
    sine[3366]=-921;
    sine[3367]=-920;
    sine[3368]=-920;
    sine[3369]=-919;
    sine[3370]=-918;
    sine[3371]=-918;
    sine[3372]=-917;
    sine[3373]=-916;
    sine[3374]=-916;
    sine[3375]=-915;
    sine[3376]=-914;
    sine[3377]=-913;
    sine[3378]=-913;
    sine[3379]=-912;
    sine[3380]=-911;
    sine[3381]=-911;
    sine[3382]=-910;
    sine[3383]=-909;
    sine[3384]=-908;
    sine[3385]=-908;
    sine[3386]=-907;
    sine[3387]=-906;
    sine[3388]=-906;
    sine[3389]=-905;
    sine[3390]=-904;
    sine[3391]=-903;
    sine[3392]=-903;
    sine[3393]=-902;
    sine[3394]=-901;
    sine[3395]=-900;
    sine[3396]=-900;
    sine[3397]=-899;
    sine[3398]=-898;
    sine[3399]=-897;
    sine[3400]=-897;
    sine[3401]=-896;
    sine[3402]=-895;
    sine[3403]=-894;
    sine[3404]=-894;
    sine[3405]=-893;
    sine[3406]=-892;
    sine[3407]=-891;
    sine[3408]=-890;
    sine[3409]=-890;
    sine[3410]=-889;
    sine[3411]=-888;
    sine[3412]=-887;
    sine[3413]=-887;
    sine[3414]=-886;
    sine[3415]=-885;
    sine[3416]=-884;
    sine[3417]=-883;
    sine[3418]=-883;
    sine[3419]=-882;
    sine[3420]=-881;
    sine[3421]=-880;
    sine[3422]=-879;
    sine[3423]=-879;
    sine[3424]=-878;
    sine[3425]=-877;
    sine[3426]=-876;
    sine[3427]=-875;
    sine[3428]=-875;
    sine[3429]=-874;
    sine[3430]=-873;
    sine[3431]=-872;
    sine[3432]=-871;
    sine[3433]=-870;
    sine[3434]=-870;
    sine[3435]=-869;
    sine[3436]=-868;
    sine[3437]=-867;
    sine[3438]=-866;
    sine[3439]=-865;
    sine[3440]=-865;
    sine[3441]=-864;
    sine[3442]=-863;
    sine[3443]=-862;
    sine[3444]=-861;
    sine[3445]=-860;
    sine[3446]=-860;
    sine[3447]=-859;
    sine[3448]=-858;
    sine[3449]=-857;
    sine[3450]=-856;
    sine[3451]=-855;
    sine[3452]=-854;
    sine[3453]=-854;
    sine[3454]=-853;
    sine[3455]=-852;
    sine[3456]=-851;
    sine[3457]=-850;
    sine[3458]=-849;
    sine[3459]=-848;
    sine[3460]=-847;
    sine[3461]=-847;
    sine[3462]=-846;
    sine[3463]=-845;
    sine[3464]=-844;
    sine[3465]=-843;
    sine[3466]=-842;
    sine[3467]=-841;
    sine[3468]=-840;
    sine[3469]=-839;
    sine[3470]=-839;
    sine[3471]=-838;
    sine[3472]=-837;
    sine[3473]=-836;
    sine[3474]=-835;
    sine[3475]=-834;
    sine[3476]=-833;
    sine[3477]=-832;
    sine[3478]=-831;
    sine[3479]=-830;
    sine[3480]=-829;
    sine[3481]=-828;
    sine[3482]=-828;
    sine[3483]=-827;
    sine[3484]=-826;
    sine[3485]=-825;
    sine[3486]=-824;
    sine[3487]=-823;
    sine[3488]=-822;
    sine[3489]=-821;
    sine[3490]=-820;
    sine[3491]=-819;
    sine[3492]=-818;
    sine[3493]=-817;
    sine[3494]=-816;
    sine[3495]=-815;
    sine[3496]=-814;
    sine[3497]=-813;
    sine[3498]=-813;
    sine[3499]=-812;
    sine[3500]=-811;
    sine[3501]=-810;
    sine[3502]=-809;
    sine[3503]=-808;
    sine[3504]=-807;
    sine[3505]=-806;
    sine[3506]=-805;
    sine[3507]=-804;
    sine[3508]=-803;
    sine[3509]=-802;
    sine[3510]=-801;
    sine[3511]=-800;
    sine[3512]=-799;
    sine[3513]=-798;
    sine[3514]=-797;
    sine[3515]=-796;
    sine[3516]=-795;
    sine[3517]=-794;
    sine[3518]=-793;
    sine[3519]=-792;
    sine[3520]=-791;
    sine[3521]=-790;
    sine[3522]=-789;
    sine[3523]=-788;
    sine[3524]=-787;
    sine[3525]=-786;
    sine[3526]=-785;
    sine[3527]=-784;
    sine[3528]=-783;
    sine[3529]=-782;
    sine[3530]=-781;
    sine[3531]=-780;
    sine[3532]=-779;
    sine[3533]=-778;
    sine[3534]=-777;
    sine[3535]=-776;
    sine[3536]=-775;
    sine[3537]=-774;
    sine[3538]=-773;
    sine[3539]=-772;
    sine[3540]=-771;
    sine[3541]=-770;
    sine[3542]=-769;
    sine[3543]=-768;
    sine[3544]=-767;
    sine[3545]=-766;
    sine[3546]=-765;
    sine[3547]=-763;
    sine[3548]=-762;
    sine[3549]=-761;
    sine[3550]=-760;
    sine[3551]=-759;
    sine[3552]=-758;
    sine[3553]=-757;
    sine[3554]=-756;
    sine[3555]=-755;
    sine[3556]=-754;
    sine[3557]=-753;
    sine[3558]=-752;
    sine[3559]=-751;
    sine[3560]=-750;
    sine[3561]=-749;
    sine[3562]=-748;
    sine[3563]=-747;
    sine[3564]=-745;
    sine[3565]=-744;
    sine[3566]=-743;
    sine[3567]=-742;
    sine[3568]=-741;
    sine[3569]=-740;
    sine[3570]=-739;
    sine[3571]=-738;
    sine[3572]=-737;
    sine[3573]=-736;
    sine[3574]=-735;
    sine[3575]=-734;
    sine[3576]=-732;
    sine[3577]=-731;
    sine[3578]=-730;
    sine[3579]=-729;
    sine[3580]=-728;
    sine[3581]=-727;
    sine[3582]=-726;
    sine[3583]=-725;
    sine[3584]=-724;
    sine[3585]=-722;
    sine[3586]=-721;
    sine[3587]=-720;
    sine[3588]=-719;
    sine[3589]=-718;
    sine[3590]=-717;
    sine[3591]=-716;
    sine[3592]=-715;
    sine[3593]=-714;
    sine[3594]=-712;
    sine[3595]=-711;
    sine[3596]=-710;
    sine[3597]=-709;
    sine[3598]=-708;
    sine[3599]=-707;
    sine[3600]=-706;
    sine[3601]=-704;
    sine[3602]=-703;
    sine[3603]=-702;
    sine[3604]=-701;
    sine[3605]=-700;
    sine[3606]=-699;
    sine[3607]=-698;
    sine[3608]=-696;
    sine[3609]=-695;
    sine[3610]=-694;
    sine[3611]=-693;
    sine[3612]=-692;
    sine[3613]=-691;
    sine[3614]=-690;
    sine[3615]=-688;
    sine[3616]=-687;
    sine[3617]=-686;
    sine[3618]=-685;
    sine[3619]=-684;
    sine[3620]=-683;
    sine[3621]=-681;
    sine[3622]=-680;
    sine[3623]=-679;
    sine[3624]=-678;
    sine[3625]=-677;
    sine[3626]=-675;
    sine[3627]=-674;
    sine[3628]=-673;
    sine[3629]=-672;
    sine[3630]=-671;
    sine[3631]=-670;
    sine[3632]=-668;
    sine[3633]=-667;
    sine[3634]=-666;
    sine[3635]=-665;
    sine[3636]=-664;
    sine[3637]=-662;
    sine[3638]=-661;
    sine[3639]=-660;
    sine[3640]=-659;
    sine[3641]=-658;
    sine[3642]=-656;
    sine[3643]=-655;
    sine[3644]=-654;
    sine[3645]=-653;
    sine[3646]=-652;
    sine[3647]=-650;
    sine[3648]=-649;
    sine[3649]=-648;
    sine[3650]=-647;
    sine[3651]=-645;
    sine[3652]=-644;
    sine[3653]=-643;
    sine[3654]=-642;
    sine[3655]=-641;
    sine[3656]=-639;
    sine[3657]=-638;
    sine[3658]=-637;
    sine[3659]=-636;
    sine[3660]=-634;
    sine[3661]=-633;
    sine[3662]=-632;
    sine[3663]=-631;
    sine[3664]=-629;
    sine[3665]=-628;
    sine[3666]=-627;
    sine[3667]=-626;
    sine[3668]=-625;
    sine[3669]=-623;
    sine[3670]=-622;
    sine[3671]=-621;
    sine[3672]=-620;
    sine[3673]=-618;
    sine[3674]=-617;
    sine[3675]=-616;
    sine[3676]=-615;
    sine[3677]=-613;
    sine[3678]=-612;
    sine[3679]=-611;
    sine[3680]=-609;
    sine[3681]=-608;
    sine[3682]=-607;
    sine[3683]=-606;
    sine[3684]=-604;
    sine[3685]=-603;
    sine[3686]=-602;
    sine[3687]=-601;
    sine[3688]=-599;
    sine[3689]=-598;
    sine[3690]=-597;
    sine[3691]=-596;
    sine[3692]=-594;
    sine[3693]=-593;
    sine[3694]=-592;
    sine[3695]=-590;
    sine[3696]=-589;
    sine[3697]=-588;
    sine[3698]=-587;
    sine[3699]=-585;
    sine[3700]=-584;
    sine[3701]=-583;
    sine[3702]=-581;
    sine[3703]=-580;
    sine[3704]=-579;
    sine[3705]=-578;
    sine[3706]=-576;
    sine[3707]=-575;
    sine[3708]=-574;
    sine[3709]=-572;
    sine[3710]=-571;
    sine[3711]=-570;
    sine[3712]=-568;
    sine[3713]=-567;
    sine[3714]=-566;
    sine[3715]=-564;
    sine[3716]=-563;
    sine[3717]=-562;
    sine[3718]=-561;
    sine[3719]=-559;
    sine[3720]=-558;
    sine[3721]=-557;
    sine[3722]=-555;
    sine[3723]=-554;
    sine[3724]=-553;
    sine[3725]=-551;
    sine[3726]=-550;
    sine[3727]=-549;
    sine[3728]=-547;
    sine[3729]=-546;
    sine[3730]=-545;
    sine[3731]=-543;
    sine[3732]=-542;
    sine[3733]=-541;
    sine[3734]=-539;
    sine[3735]=-538;
    sine[3736]=-537;
    sine[3737]=-535;
    sine[3738]=-534;
    sine[3739]=-533;
    sine[3740]=-531;
    sine[3741]=-530;
    sine[3742]=-529;
    sine[3743]=-527;
    sine[3744]=-526;
    sine[3745]=-525;
    sine[3746]=-523;
    sine[3747]=-522;
    sine[3748]=-521;
    sine[3749]=-519;
    sine[3750]=-518;
    sine[3751]=-516;
    sine[3752]=-515;
    sine[3753]=-514;
    sine[3754]=-512;
    sine[3755]=-511;
    sine[3756]=-510;
    sine[3757]=-508;
    sine[3758]=-507;
    sine[3759]=-506;
    sine[3760]=-504;
    sine[3761]=-503;
    sine[3762]=-501;
    sine[3763]=-500;
    sine[3764]=-499;
    sine[3765]=-497;
    sine[3766]=-496;
    sine[3767]=-495;
    sine[3768]=-493;
    sine[3769]=-492;
    sine[3770]=-491;
    sine[3771]=-489;
    sine[3772]=-488;
    sine[3773]=-486;
    sine[3774]=-485;
    sine[3775]=-484;
    sine[3776]=-482;
    sine[3777]=-481;
    sine[3778]=-479;
    sine[3779]=-478;
    sine[3780]=-477;
    sine[3781]=-475;
    sine[3782]=-474;
    sine[3783]=-472;
    sine[3784]=-471;
    sine[3785]=-470;
    sine[3786]=-468;
    sine[3787]=-467;
    sine[3788]=-466;
    sine[3789]=-464;
    sine[3790]=-463;
    sine[3791]=-461;
    sine[3792]=-460;
    sine[3793]=-458;
    sine[3794]=-457;
    sine[3795]=-456;
    sine[3796]=-454;
    sine[3797]=-453;
    sine[3798]=-451;
    sine[3799]=-450;
    sine[3800]=-449;
    sine[3801]=-447;
    sine[3802]=-446;
    sine[3803]=-444;
    sine[3804]=-443;
    sine[3805]=-442;
    sine[3806]=-440;
    sine[3807]=-439;
    sine[3808]=-437;
    sine[3809]=-436;
    sine[3810]=-434;
    sine[3811]=-433;
    sine[3812]=-432;
    sine[3813]=-430;
    sine[3814]=-429;
    sine[3815]=-427;
    sine[3816]=-426;
    sine[3817]=-424;
    sine[3818]=-423;
    sine[3819]=-422;
    sine[3820]=-420;
    sine[3821]=-419;
    sine[3822]=-417;
    sine[3823]=-416;
    sine[3824]=-414;
    sine[3825]=-413;
    sine[3826]=-412;
    sine[3827]=-410;
    sine[3828]=-409;
    sine[3829]=-407;
    sine[3830]=-406;
    sine[3831]=-404;
    sine[3832]=-403;
    sine[3833]=-402;
    sine[3834]=-400;
    sine[3835]=-399;
    sine[3836]=-397;
    sine[3837]=-396;
    sine[3838]=-394;
    sine[3839]=-393;
    sine[3840]=-391;
    sine[3841]=-390;
    sine[3842]=-388;
    sine[3843]=-387;
    sine[3844]=-386;
    sine[3845]=-384;
    sine[3846]=-383;
    sine[3847]=-381;
    sine[3848]=-380;
    sine[3849]=-378;
    sine[3850]=-377;
    sine[3851]=-375;
    sine[3852]=-374;
    sine[3853]=-372;
    sine[3854]=-371;
    sine[3855]=-369;
    sine[3856]=-368;
    sine[3857]=-367;
    sine[3858]=-365;
    sine[3859]=-364;
    sine[3860]=-362;
    sine[3861]=-361;
    sine[3862]=-359;
    sine[3863]=-358;
    sine[3864]=-356;
    sine[3865]=-355;
    sine[3866]=-353;
    sine[3867]=-352;
    sine[3868]=-350;
    sine[3869]=-349;
    sine[3870]=-347;
    sine[3871]=-346;
    sine[3872]=-344;
    sine[3873]=-343;
    sine[3874]=-342;
    sine[3875]=-340;
    sine[3876]=-339;
    sine[3877]=-337;
    sine[3878]=-336;
    sine[3879]=-334;
    sine[3880]=-333;
    sine[3881]=-331;
    sine[3882]=-330;
    sine[3883]=-328;
    sine[3884]=-327;
    sine[3885]=-325;
    sine[3886]=-324;
    sine[3887]=-322;
    sine[3888]=-321;
    sine[3889]=-319;
    sine[3890]=-318;
    sine[3891]=-316;
    sine[3892]=-315;
    sine[3893]=-313;
    sine[3894]=-312;
    sine[3895]=-310;
    sine[3896]=-309;
    sine[3897]=-307;
    sine[3898]=-306;
    sine[3899]=-304;
    sine[3900]=-303;
    sine[3901]=-301;
    sine[3902]=-300;
    sine[3903]=-298;
    sine[3904]=-297;
    sine[3905]=-295;
    sine[3906]=-294;
    sine[3907]=-292;
    sine[3908]=-291;
    sine[3909]=-289;
    sine[3910]=-288;
    sine[3911]=-286;
    sine[3912]=-285;
    sine[3913]=-283;
    sine[3914]=-282;
    sine[3915]=-280;
    sine[3916]=-279;
    sine[3917]=-277;
    sine[3918]=-276;
    sine[3919]=-274;
    sine[3920]=-273;
    sine[3921]=-271;
    sine[3922]=-270;
    sine[3923]=-268;
    sine[3924]=-267;
    sine[3925]=-265;
    sine[3926]=-264;
    sine[3927]=-262;
    sine[3928]=-260;
    sine[3929]=-259;
    sine[3930]=-257;
    sine[3931]=-256;
    sine[3932]=-254;
    sine[3933]=-253;
    sine[3934]=-251;
    sine[3935]=-250;
    sine[3936]=-248;
    sine[3937]=-247;
    sine[3938]=-245;
    sine[3939]=-244;
    sine[3940]=-242;
    sine[3941]=-241;
    sine[3942]=-239;
    sine[3943]=-238;
    sine[3944]=-236;
    sine[3945]=-235;
    sine[3946]=-233;
    sine[3947]=-232;
    sine[3948]=-230;
    sine[3949]=-228;
    sine[3950]=-227;
    sine[3951]=-225;
    sine[3952]=-224;
    sine[3953]=-222;
    sine[3954]=-221;
    sine[3955]=-219;
    sine[3956]=-218;
    sine[3957]=-216;
    sine[3958]=-215;
    sine[3959]=-213;
    sine[3960]=-212;
    sine[3961]=-210;
    sine[3962]=-209;
    sine[3963]=-207;
    sine[3964]=-205;
    sine[3965]=-204;
    sine[3966]=-202;
    sine[3967]=-201;
    sine[3968]=-199;
    sine[3969]=-198;
    sine[3970]=-196;
    sine[3971]=-195;
    sine[3972]=-193;
    sine[3973]=-192;
    sine[3974]=-190;
    sine[3975]=-188;
    sine[3976]=-187;
    sine[3977]=-185;
    sine[3978]=-184;
    sine[3979]=-182;
    sine[3980]=-181;
    sine[3981]=-179;
    sine[3982]=-178;
    sine[3983]=-176;
    sine[3984]=-175;
    sine[3985]=-173;
    sine[3986]=-171;
    sine[3987]=-170;
    sine[3988]=-168;
    sine[3989]=-167;
    sine[3990]=-165;
    sine[3991]=-164;
    sine[3992]=-162;
    sine[3993]=-161;
    sine[3994]=-159;
    sine[3995]=-158;
    sine[3996]=-156;
    sine[3997]=-154;
    sine[3998]=-153;
    sine[3999]=-151;
    sine[4000]=-150;
    sine[4001]=-148;
    sine[4002]=-147;
    sine[4003]=-145;
    sine[4004]=-144;
    sine[4005]=-142;
    sine[4006]=-140;
    sine[4007]=-139;
    sine[4008]=-137;
    sine[4009]=-136;
    sine[4010]=-134;
    sine[4011]=-133;
    sine[4012]=-131;
    sine[4013]=-130;
    sine[4014]=-128;
    sine[4015]=-126;
    sine[4016]=-125;
    sine[4017]=-123;
    sine[4018]=-122;
    sine[4019]=-120;
    sine[4020]=-119;
    sine[4021]=-117;
    sine[4022]=-115;
    sine[4023]=-114;
    sine[4024]=-112;
    sine[4025]=-111;
    sine[4026]=-109;
    sine[4027]=-108;
    sine[4028]=-106;
    sine[4029]=-105;
    sine[4030]=-103;
    sine[4031]=-101;
    sine[4032]=-100;
    sine[4033]=-98;
    sine[4034]=-97;
    sine[4035]=-95;
    sine[4036]=-94;
    sine[4037]=-92;
    sine[4038]=-90;
    sine[4039]=-89;
    sine[4040]=-87;
    sine[4041]=-86;
    sine[4042]=-84;
    sine[4043]=-83;
    sine[4044]=-81;
    sine[4045]=-80;
    sine[4046]=-78;
    sine[4047]=-76;
    sine[4048]=-75;
    sine[4049]=-73;
    sine[4050]=-72;
    sine[4051]=-70;
    sine[4052]=-69;
    sine[4053]=-67;
    sine[4054]=-65;
    sine[4055]=-64;
    sine[4056]=-62;
    sine[4057]=-61;
    sine[4058]=-59;
    sine[4059]=-58;
    sine[4060]=-56;
    sine[4061]=-54;
    sine[4062]=-53;
    sine[4063]=-51;
    sine[4064]=-50;
    sine[4065]=-48;
    sine[4066]=-47;
    sine[4067]=-45;
    sine[4068]=-43;
    sine[4069]=-42;
    sine[4070]=-40;
    sine[4071]=-39;
    sine[4072]=-37;
    sine[4073]=-36;
    sine[4074]=-34;
    sine[4075]=-32;
    sine[4076]=-31;
    sine[4077]=-29;
    sine[4078]=-28;
    sine[4079]=-26;
    sine[4080]=-25;
    sine[4081]=-23;
    sine[4082]=-21;
    sine[4083]=-20;
    sine[4084]=-18;
    sine[4085]=-17;
    sine[4086]=-15;
    sine[4087]=-14;
    sine[4088]=-12;
    sine[4089]=-10;
    sine[4090]=-9;
    sine[4091]=-7;
    sine[4092]=-6;
    sine[4093]=-4;
    sine[4094]=-3;
    sine[4095]=-1;
end 

// ROM Logic
always @(posedge clock) begin 
    sin_out = sine[phase_in];
end

endmodule
